`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rDtsobuIlJULUYu2aNgvf2+P/kC0uC0I8zNOVL62Qqf7G/18fCRI5auEOITsj2Vr2hFVGFYLKhL1
SBQ5U22Awg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SGEzlu7dxmwGcYphI3L3R2NRZ6L+FpSO3J2xi6Mws/kD1bZST5DxeQOTAyp4ts0eGq+PMTwSfIDW
NbyYrxB4EJ4zg1aQclvACH6sKrrwepJMyFk1Ea7k7A/uL45k8A0PGAowu/IaOKbL/lTSd2xnCS1v
vPYLrQGgoeuA4yYfMK8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
17dL3KnCEjrp1c77oZ+kJjbT5UTwnArewt71zQkDttWfJXBWEC3ySJknSnXnb/GVJjMnfhyS3OW3
A9VxVckuAEITGYg/IQeltik31UvB6uLZoaznsd2xa1YMNnq5M6FMeYN9Wx+u7LXZyPemVcEtVSe9
atXZdMbPoeKVXOFX6RJz1OwS2JwgZAWXR7Izo8KAALCxUvUbFCfR9TSlLBGzeXoZd+QYkm+AJLxb
WN3zWfErRUVg+04Vh0q4S475PHza4aXAZTQkWQnnBJxFDVmS+4xYDKBmA32T4oh4h6EGQS/4jS7h
5hh7IwZFX4oQNbeeCzYCS8f6SGIOAzcyHTyNTw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e5JKyDNFpXuNXCDfnpCh7rmH5mRdgNH1dZ0a9LcRKLWWKj9HZqG7BktAzETST+yrbjKsxSkAjvQJ
Eq/6quIaKXU25Yj+X0Q52ot2mOnJRclQyzQGKJsRxFnp8NqpzczeP6oO6zxH9Ln6aGpowWFKrqRd
D5DIB4ALLdk18yWVveYvaj9n5V8WC3EoHabKWhDT5dt0bB7+DBoXq0eqaX3ycEnaxPz3gs7/ZfQ+
DV4VBrHzkvN2kUS+qhYH4ZFbom3yCZXg5z6/GuT7SaJEWNj5ToG2vtIIA8wwoFhP5oJ24eDxOtaD
MPOeoDU7PZAK9984F/oHazsPf84qkVNFYlAd0w==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Dl6TX/MFTTiCU3BWAqjWdiuyUZXOoy8N6F5PlMEFJuePUXWN2gkmJp2ebA1q4s7wa7UHtwZsfkPO
RrkRV4iB2IKX7MCuuEvcDAOFPfPOI+sgO9GNmPBW2mU1hZneZ7gOx7mrYIGvNc+3jp6guuY16+b0
un31GhBVR/+DDQfhjLrvCPOdQvxTkVU8j4LNJN3HuZQZJ4AMxn2fE5WATeEBScZylAMnOg0D52Bz
eeQlc14lPvYx6FtZNaN9k+SJ/eveH18WXqE+D8G5pyb2siBdPdpP9qhl5oqSDqbVuRxGKoVDgk98
9Wg3zXYtlXEle3vvXqzk56LlfCtRPAsUzOXWVQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hBro+TIeqRMnluKdDuU70qnCxZmKu2s3BPsWG+NVU9zNJLwotJjtFNmwpTEHCIuxcgEV6tmn3zSb
MY9yfG4u6TWepZiGCbhv14vPsWlYpM1MOb6Lqc2hefEwGQf6eNebcZUBZE21KPnx90MDbWaE3Kj3
ZknDvUA+BXhHYk8ldZw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c0W/m/n78VhNb0tgozbh5krwuQUnCXfaDhHCw6DMykQ5RbndCvxewQ3Hjd2ikcXg25ApN2vQ/0s7
tf4xFiemrmKCtP6kFnS8+eh01nuWl8AMWMiCypQ+GbeJyQR6z3f45WDIRYlHYcSjinUqMy+GYTSL
ITl0J2djXYMZRyPxFkFR05s3YQAnYCqJmP6TTED6FllxQ1ZFVMQAHIC140Kv3MKHiYjAIuX8gtdn
Q3H59eKT+ORXIhTwMo8AVQ3xs/nr8yLqXlM+6yWj3UPiHOaJlZSkkdES/w3f6CWGbee+e7u8+KVB
gLsI1DI1BxNYO7mBBW+fi87bVHkhcX5Y8snpBw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432800)
`protect data_block
m+uscW0pEk6oS7BkdE/SVZuvg4K7NYZMg+4o6y23t7TV6W+U1JZ9E8LK2ZKTubAm7jNMMw6MRhD7
OPgJoi2opg+JMW0eb7nsJzBoUV0gdofj7YnzsruRhOnb7i8ni1k+qmVbBv4KKecpeD1BPyoeDhMp
6gSveqzJgKVs5sO8jYNRHHgsbQKMYAulWSEOuEMHNv19/nNBTUkC7ow8bxCt7sixyWCkIz1CvbtT
1e3uWBEYI+53EQ8d8Z7xeLxYXYYbOft3vJvYoDu3JaagqfOvN9BQffIUFmemdEsZWosJL1/JM7+Q
LqeC7gaPe5l40ML/zW06Jk+I300rPr4WaDK25ayiDCUJdyTU2/Uwrn3meqw/tPa5E6wDR3Y1mLlC
WakZ4kSkPppjbroGaQm479+wGeAL3A2STWIgdULkEP//RHCzNmkFv5Ea3l5OnQVFnIj9XeZ6Or0l
UGP8LwxI0nMf7gGC5BKuojThVPmiNqKKGjVtG40StbFtNsDBEQZ0Ke1XpertcDazwlsVzAkkcG7f
C5KBfIQobHABjkVSe8lUO7kO7ANr/jXnQhykfZJyoDs79tX22FKoMXrDrBosFXlrTFegmZbdDDmb
4eKh+vyuddE8KRJPK8SvNnJKsEWm7W4UOKq1Mi0ruQ94rYMj/S5wQOJaDrsJm0NrEa1z3iNAOWb+
mAFZ9ak83bYMxpoCW1sM91WmEEIVqb9V5j/4nCv3KmYjBAe3ApKK4P1Cra8xVg3gOY9UxBPfCi/9
FyUkMaJLKeapdbC+MVHX6U7wWcHkZAFFwnfJlohJwkJ2Vg2MPCPi2sWSZ1lDzTr/djFVOJw7odFw
zvmPhNuRg4+2MWss7MpC1SwQooU85CXDpCZL5UV75LRL/mD10wsrmGbBSosm2+E9xOIBzDteg96L
gvSAgkjL4VMfn8LMbYG6b1x6am+wVYsSB50H7wt00xHMTW7n2dag7322XXH5YvZL2YSprkB/5tpd
fHxDY5ckJPYwMui6MDtSzT525EGwK8tQe2cJFVIzHEm45fU6ZVeTCMUdfuD0sPFcUh+B9T4Xgeok
ay4Ix4mAkWYEz/skUd6jXQVTnoNIn501nLKm8tMZ8IbQY665sUfamQZUiuXgtu/eTPa2hKaxHwwL
pPZa20E01S/1LhI4qSxW2KsUXG9EVRRLY4oiMb+73obiVL9/rUTA2xQzzsuM0ZUybf8vdVIOb/Vi
lUbAhFFyzBL9aCoTPqX/qiHTiNkkTjZNktGxxf8gUr2P5IM+oOpRP9xLFDnXAne03U6iDco5eDp7
LBF389utRjtO3uZ/iMi1jTPkZXnI7Nyw4z545FwKBm4PUl0wEHavrux2BN362G0U8GglL3Effv/a
P+EKZ2Y+CdVSunyGiJtgkO5Pgzoi6uswaKqSiRbUKAZBns+n6wnkfKWSNU5aAA3xUW2PQK44Rxjz
amde4u+mcZ3pGaOA4AAg1HNvEVNZ9uAIbJNlodgJSzFKvu08/fqQHIwJprsLYvcMYAIsw3XycvKM
i+emhsMe9j+tMbB/bWGu6qhQ8ZnCOZNrY5pSC9wehPOMqELcNgwwR7t+S7u61lVrw2gH70eIQjpZ
sAlFkvTkMKu2m8YZL7KunWylOGXa0lPwwwKh/VQ2TqQaotSyDIDN6qXycZ3puYd8EQPL8Q+lhU8T
5PVkUO6JBhoHvFbx+ZjE45lVERYmIfo82tJ2ClBtJDvbG9CNGCnVyXIOxoxTQDQM1vTAODWQppP6
3eTZo01enoTnwaGswiYZOB7nxZ0S6v1HiB9qCAPY8quG9p2WG5wZhJAFJZSrxHJ/Nd10jrVros5a
Ac2USP2P1j65CgTr6bppjbu+0g8NFOB607+rtiEIiIwQR5Sr9CTW/C/UKdBegjj/SSuCXsX8jXUd
OGeW38Eg1QhMhcGgFCRnUf9U091jqvTf80oMDFMmlfqeDJ3PaI8eDiqg2Q/8Xzi0tkO+kEzt11gh
7+tC93Dhg5Zeh7CPjRtRCxwrzgEyCF2AP50cFkGyF6bj7D/2BmwK8eoTIxYAZGv9i/dnMbrwoOlk
jGq5afXd50ErqI7lp3FoL4hAZ0sSOhKuX2Ebef9s+kv7arBEYqpRQZkQWznyJkIdOJIKEYtsuGT0
s08NEQV/we7AobTSdiHZ4EOZgJRCCi2JUlv/A156gNAs5BCd16Sah0jBvk6rF6BH6uGp6c4FAuCM
T1GcmSekGZPKjFc+rOfjFDITqj081VbqYBBBd3eem3w9m+8CPvqrHcD5SiZ8Vm4aHkuReHsE25kk
ctC6rBOqES2eWKcsu9EN9JpRo+0ainLgHPgxnVUrA6XUrq2x1KJ/uLbsVX/vJX3L4lHfBiN2wJ8v
kQG8qHQhWVvmV2KSuo1nIZJkuPtyj3JntY4o1QPgaRstO9+qn7VOvaGyoBw3ahO/GZklQRcN7ygr
IARzmZQGiwC7LKBp6f47qBNFthEQ7/Ut13U1vG8O00TkRqqAAxck/aKje1d3yDa3fDJf5PkykUeo
2l9ltWK4Rb9rkFftYYBMMyKjt/Pl+/nYfbYD9MIkN0ssKJZptPDEoLZAHZd+lTTRYCbUnG6h0bSD
w58z+JcpnGyL92UFIWg+TM9/0/ed2GzGPolVvDAK/nzkQ1Vsm3JmB+U8MKpje+brRXZDShDKldK1
3oTT1bgIzCVPHq6JXI8LSHt3w2z/Pl3UUq9eOHGXmAgGbbyNjAuJNe7Y2ClMY/hOB46apyd0nLBj
aOFQX4iaWHpGEeXtqNk1HAHyTh2Vu7/OVxEIHC6C3YyV83t+mdupE+YcveRGKByPSpuGzFRXpPP7
kMCNlJPmp5pslI0PFSRy22DEoywr30L5SaDw2o2A/mbR3vPki5ucYEnriK+MWBBAx8Q+BVfqSQln
azkOxGw8ZPDggCkfVkQLXzBzCXm05X/z+apUk931ELLjCfgiqL5O7YIIrh1A2uHVgFT79PifH/rm
TisO15hZ25NyXA3rdwxLcE2/IPpuCXl7arY3sFxEF2bhxeLB22QhblJGYDKl03Dq6YjtUAfXLrKD
29XYXh55W/PG8opvmLDV+WiqcIJ6ZWpUtuL1q4QyIqAzudwkA+ZA17Q2+wWQXZnPS8w/pc4gy6Ll
mJWN7KpTfzXFWedKda1uCMDhBpAiEfbKSPCv/I+5DHuP/HN10tI0dhDybXIfouTpppiqIIWGBD8J
ZkuFWjSZL6pKkqXoHZpLyYyx0GE9LSieqtH8gmqcS4YaR/v2macz5If8w4F+2NNBmV80MBu3co2V
DONvoHOpH7U0PWc8aWMzrDlIAjPOaZKnRZDUzdMaBPkaC77uE0v4lA36XQwunu/3wmeQv0AJ+KGf
PHJArLlY/hGN/tmuBLATukdkLCff4BjN7fCcVfBnWn0LFaN/mZd8aMq+J7Jd+3vW9q4pNsrER0ky
b3rKx0FwEC4nVcou7+FLxYJlPYRr9BNHQwE0nbhcCM5hjQF0EAC8N0D5Hb8cfUx1LndP6L0cpoHb
p1cATL1Yb2FazMyXyasaw44nHEkhH3Umq0xyV/dN4+3hNczf1a21g6bwxpWerkbwCTZlpcUhRbPG
LmcW9+hCCwGq3L1r7lyjEVTZ5DsaEPMHRmXOvdzrWHMivAvXBhez+IdQ+uw7KufA575ayj70Bm0U
1YwdNOr0VpeUVF7zL5kJBCRoGbOOev/YZfYyqITOVrUD+Ij1GJq1yHLHkk17vz3Uq0+K+ajjzOyF
5HmcCIf8O1sib2Zuwo+qBQ+IIuUVbDkpbGLYC4DaDpW/A940O4STjbdiqtHcODw1wGXmrgg7TpUa
16YKFLE8oHrlrGrb9esOmFfGWYt5YDmJ2C/gDTg0gDGapfomuHcv56I7sGX6ng3jFyvOvb2jS39c
AyfnIt1pk2wjZZ7GhCZi3G8tR6gjnBIWgCwxw5ZtjCGv85iQdQmfPi27F7dOT/zEMHpeBv+YRd7A
rvnH14WhOlZqEtmxzrHZjf/26qbY2tbk1bXGM7rVM6yfaW23DvhZ2iRJblkAwRQeFq5PR639ult8
z/66RWqiz9YsXbPSj+Z/VJaLwCGHQfJbRr5VxLtZda5ZfKIral2Z2MWUYSlVv/I++N2JGdsYcX9c
/OEuwN0MgumlDUrWEAZxbnnU/Bbbq+TGEBGk6tvfcPvNYBjOLhacKuCm9gGg0PShi4jaKqvC4h7k
6WyVUZKU8KArD2kUDvygHLgoxYqpTuFEZoCo26R7nbjzGmm0Zpgpk196dJbaeHpk4GfZ9BSlI9Nk
hRA632mSsGp8Vqz3uydDy/QmBfWubHBdKzSvXU1O4CuOpiRY2CJrTsgwTqHVY73Xc7Mq7InuMBIw
x1PeN9JGxBPid+OE0DMhPH5IhIVlXWUmI4I9awcr+3MaS1gQ2iRQ56IRNZO/MtwUPilL9Gckwrtz
lgSz8aBFj3dvRYJiKRzFyh/Bd2fmA3tDGM9y/BP3tBKiLmb3ziiAlDjrqmBrc/CYasOAsSh87diC
U5kG7ny56BCwWs8J3KPzwCfFDN0L9NTfoW9YNgxFDr76uE/2tzJgkRPC3OHfcy8Axxk4tnrkyiXn
gvyA5ZjYveElMPNjpWKeW2HzWoibbnygyK+yJYKUyOYgZJgK9SyVJljFkq/8HkJAgj0Xt8KiRZER
yO3QHmuX9eq3jPOY3qGHJkSbMbx3/phNHJCpxYceGbX26b2b2jLvLrXqBz0wnXSNR8cZRDUwD92b
zFgIi1rrfrnA8oUmLMwbIDmLKw4GfZRqox02IdIZclaUOdXDlX3SIRKolmPCWdJto89ebYNcn/I3
yscTgsrUHoMQrYmw6k9gg6AKD0vr+e2C1ZhfU082L4xP3Pcuf9tRPRBO2bi/zzmJJzdQyJdM1iQy
Sy4fLnb2aRpJUnt3VNTcpj1xu7TSOyYD2qJ4+v7uP/mZTFfxrF4Qipe4sUSeTycLxNkHxo/GV4iC
Hf5WTVbxJVFIGesnFZV6jTER+eYPPrkz3ftPi0GxxN6z1jmRluQDpHcDZq8VukOs4qmDEPuihbhd
SbXg2m+9QECciEtPKsFsu4mGgnN7n1bWOfT00pLh6MF+/3AKcMWNT+KL6yNVXYnEnhguZ70RsxvW
pRSdGWd2Z6jO+wx5LSotrlTWxTbFNY7EBG737gGF0vg6SazNam16paQVyfGTyJei7o+NXvNF2EwR
RIUkCf/4b3bC2Wgc7DwJ4zA5e0IFGwgAu8fer8lF+G0whSmHWKnVfr2IMfSks+y+9ojYx159hTor
VkxOHvRplZtpNYJ0PgD2cwuYXynuKs2oimsSywom6gW8cLieLxiaREYuMHHfR1olBR8FRg+6TxEe
iUDIxsyEI7bUlvqD2z1PkmpG8rRx0yOIBDCeSNhh6UjY2aeQBznHiXRVu8CPm2Jh/ZgJGWkupdP+
PcqNrQjWLqkRmUWUm2naJHO1iFnZCK3oTqMrNLOlhVPlCpo6OL2ldRhgJEXrH8vN45P7gQKTgE+Z
WEi6eeCLthMo9tYbPuuIqXyXdz8YPyMlFYpci09Y+pyKCL93l5XvcZYOzdeI44gGy3oCehIk4RrA
RL4dpGNkjcdyaqB5JRzeDRCi1URIQHtAvaoTzAwPunxwSpCIwcgPEq98rmFCA7MQJZAMzRulcuWo
9oTUaBrcS9zaRu3LKpEog4e86JIBDnRr1I7Rpc7+0v8DRysHtzlhwQxnF3WOHCA+PCqljfMe6VWz
svAVShm+k9E0pX7JCMCGSY8Lb69UCDznktsDMX+4IeOmeExrboBZWGvUxmgjHb97RKSLXhF1rE96
zGIQKwUyPlsq11sw889pT8Oqw20HaeVEORAftOi00b2HuXrSr7tIo6iPhUhcLzUoaqWGpxoab4qO
9RgAm8dOq8zalC6+l9Ye9qEhKlI/Esyx/HA9FJCsC796QFBF3ZArwEL33OC4xnA6EKAX3pVqqHWM
c+uBbm2g67wN3dOCmLNUWLuYhwMWa50IeDyqbsVGoUj/QE3Wa3LKFKHWhaXpGmXBCJ/kkdEJoffx
aOcCBY/EC6iiEARkMpn+RMKk8OrMf5q0GKJdZ02D+PuhEJ4NK/zReBVIQOeXzGGYsOpD6tkwjK+d
oNegL6hbW6eD/01+I3JbQ9ZhXiGohENkyxiNdgKDwrc+CWLR+FVqFej7BG1yK5G/T8YleHRcOlap
B78vxNwGLhcBkHGzlxYMdLIVaIylXWvBTV5OCdQJVsEF3ua2n21DAxKEsmlaEuzz+gHVDE/maFZb
RFV4CQz9MeKKnHho0pfEqnvC6J5YexzRGxSK81pgGvHV/de701iYOhnVRItxRTBPi3q+Nivpccy9
4J6vGLL9H3BL7BjN01cFH8EKGprmcVd2KRpnX9mQU4AJPa242U6VCC0eVPhrg1ncZnwyq0luH8VQ
D7tlI9SgIFVvAGwrDPAI2FCBPIHrH9gs7/hYxycrU0PWcZNRBdFdEIy+uD87UVAI2FGCdIoGjdtH
IBSJqOzAeDAO03f5N0W7H+jzhvgNbAI+9sMhXTbyLZ84IE8LpfVAviqMvFsl5B+FCJWp2rejcQxY
OjL3RW0YyXr0DKnsrG+lTMB7Y3z1qnAHKPOmpCwLiNW+dyHYffjNaq4XIv61XcpuVcn5PZXTfMPN
rOT8CeXoMp6DzB8CrzjRCmLcKwdrKWzzf0E3j6pPt/i1spD4YgxvdBINqv/prqvEWckzDhTxfVJy
eqRc2X/DVulRMdChnmDFDts9kX9x38Nh7OKKVAow4r+HVdAPi1hdZA1gUgnO+/PWPdtAF94YETzQ
yRsFOJqEfZpp4MIOiYIMO42KgAcySqC/5sSlOdh0RhgqM8I1DZwIrH26oCh0rQQwOm93Cr2mpOrY
q9q+rMFOrbyQCowzy0t5Z0+07HeH1YESTq3Z3eGXyDOZUbe8hmqwtYO8ErzgRabG6AT3wPwxkbtP
TWcmCH3ykVm6NGxAhpkFATDKntlD8EqmMgHgNF3stuD8WmURc29M0LPfsMpHw7eZ8h0goD2BdRh+
F+pyWk7ZzKf8uJSS887vdNjr8hfsNNsLYnAfhQHRXQWbHtjmUvlodD/495b2B3MTQv63rl/6PhuR
Wm27laOzxfB9Vq1EbK2x2Z4m5RFcscCJ/h1GjnOhZo+fTfjvYF/JW3v0WkXnIJp54F92oXELdMCS
hBQiVvUwvIdSVexQ3H2BJrnbS7TjqikuP8OZRcKtQnkYr4NfZof/tfeFDRL7tCkMquTT6sUI3ZNO
Uh/BKm4qWV7hClYrC8Jt5wBW1AJOFfV/hZVQDfroqXk3weYZiEQqVn1sio+qGIXHaAs4DPwc1UJt
aYFl9dHx0QC3CjIrPdqrTwFcHOa6pXAgrsU9BuYIraww4iVYRCZD79Yz9rYV33AeaZxFcgSFu+kd
7pRRmHTiIOeg5i1UfvrrCqHUXV2JOpi50n+V8n4d4wCDUIx7rLSMTK8oUAPis9HfroD1ptVKancv
6EM3X3a3PhFHjJt8/nbO20YZiprMoM4kYB3ntNBLI68TOHUuAbld+T9KQdvtm2eWVCceyQO3fx5V
uoJ2b34aQVFzXPlv1FeeTdIepQuxVTX7RJBrOhTlwD4cYDdJ5sdoFJ5YbyfHoMbhk8ZzFgaH8fZw
NHJhxxGZfrxnDMizoG9jv0/KgM8FjYIBnrKhqhYFXCuBlMtwsNFZqakINd53aayzYlzvpHVqASLM
1hqVPdxz34SM0Cc7tIQLEbELxJB9+vd72tC/YHOWJNHCsXpVBhU9BrHqVuFVjY2/NOo87Y4voC8I
OJNEjnvHrFZf5L2UW1GIb1xBWFPzyzo89S1UynW7kQxLxzDlku2Bt1K7Ny24YPnewKmX3XwL06bB
amZaiHsYvFUSxlC4xbwIzgSp+2FuKGFewI7AjCSnBFsOhwX2yhmIVudaSfiYWtrnRIpUFgLM8ieE
6dILFDPW7z7Hcg6hMT3rOc5u7QVqhrmvQAT40hI4arRjXMNxWNbl0EZ9ZM2rZiZjaOIHGnYTLDAq
e+ldpi6zV/yXtN/Os1BXTI8OenuSNJW6NNSPms4zfahaN6E0Kd39+0zShMKfrYKkJ+zv88+4g+K0
QqUxSBfEZ/qjw7z5aaoTAVoqRkxbibyMYFwFMm6kSysIWMI2URQciN5NXcQaG38Sr3m0KUU2TrNR
hQRdnC+wZsW0t8Y5fvQLYE+aAR1/FxvynKTSrESfzSzXI2rQaJev78yR5Ol8d83f9T7Cg8wW/8sb
RssEbdXhQRiu49Nqvoj+D+ul7krRhvOFyHUa7JqWEmsAqsOAnYLfAFNNPW0UMKX96g1qonMsomuP
mCNtvdO9MPreu+JI4f8GpETUKYH0e2T0F0n3mAcAtl3mu03qDvWXClWEc50MDBogmBprKSrZJ704
rxV62H4Eun2NO0xQA/OQHwWu2B2ZfgdtI7A0u88lVEexWWKJDd0ZSN6WgXmKRW1WNSp0dM3CE+Hw
Ujxp+muXfjerogJm+cRw15/XVIlAcQ71B3YrKc8hc7u28zpFk13FwlEvt/46QESmtwG6hI1i5dYa
AYt09v6AyoEwp54AcgUjV3CgYsvXDAzt3D+lLSl38OLugtJR22+/V6/Jhm5O6U6DuriclKf+Dazi
thzSO51b81VTOYjbJ0Zh7h7iZbCzA6AREKmH9XHrt2pDV5e1rxCuteXR90z1/BW+Z0MHsB5kRitG
FHpw2szLJB7bxm/AMmz0CXeVA42J0k4g9iq/RyDu3dsFVB8PmxZ9q8xNmX2y7jQnP/hHVA1YzYJf
FKPHVSuglGQ00bd67mLiuGquMsZp29/5jTZh7zFnilzGQTHQp7pvtvMBdt0CJER4IecCI23I7n22
q6etFdDzCurEiCNUHqnBkdVIqr3TqKghbPQSU9wP2ecaHPUMIQ621pnMLzmvWO95fnQj0BkPhizQ
wHvBIZAei6wwEYGSbDW2UfVsFMx5ShBDwUcvh8eFtg3VQPswBaJd1PmvL7zDMpnck+Bzsd9gS8nZ
6eghV7ziOckhmEumEM15Iy3M6cQRQm1UlqYGHGAwU563U+vDVTPDDdHkSe5gbXtYzBYqGYhV4I+3
p/c4xCuUuI3npHw+kuNVs7gBdXYz3BK7VJvFLV1Cr6kYumq0Oi0YSgs4XEcT2XuSPiFIhLh8R8+H
qb64t4OgysbSkf0igZTuzLbj2LtRiLqx46+2SUhYPo3FjR8gH77D+77o53Gp3KD5KRogx5+mGZfv
GaAEtgwJVrq2pA+xzXiKLonZWGfiRn+xkGwsi4EyRUSlVR2MDGkpuQNCqmRGnztTROM/QcKtgEf9
16WBJDanz6yAKQGZ/N/tyVwnEGrXEZ/blsoG680nmPMm5Fm58TszGcqa82cCYvXsSC2yG+A8GxEW
zUK+A6JZ8g+81tSn9wOr2QU+Xx4RQXmRO212oLvKcNzOSZo7jSBDtBeJsnfA2X5dTKlhbXaquSQT
lBTqHEizXAmlZwyR4NGX7hShEAOLceJ3eEx04NxKNu2ILNFIlEXKr/wkhnppIZxNpYj3p5i7qsMG
ZkugxDmAQGbLxzdSk/wNxv5QpekbdkIzDNrObj104FcchPtLYcvacTge7a+ITKdJ8oUhr7BiQD9t
gZ9NKlQ8LH47tSHvOq/HG2h9Ycp/PeOhFQ8Xe7tEQ5gUYCgpt3x79Zis/W5T60Skkh2KzvuFBL3i
r5op3T1+Yiyd9mR2dHEUVj4z+jepOI68JgJWgBN9Ku+1r8L5d1cDCAOW/P+2AKIJbOOnoZoul0MM
L7ZBXCdzS9dmcIdthNERI9Qk82d3ScMP4HyOMv7a6nQ039YHdfsWwfd6G3yk6ofbumpkEO7MDOo4
sAFcNZXnnAQwkxA9fdK+5cZtIuUzKxvgVA7Z7LGZMbrwDwc5gyA2mO0vPEGDH7cAo8u1NGkuJYM0
Ta52qsE3Vi3IjHJdq+3nsIHtn/9i2G9CEKIVVRWnuUWdm5QXc8C7YuNzxdd7UD8XQFjp6MViWs6E
QgCf+vlPqN30YuOgFvLocCpbsrSgWZCwPoPmfiGvEfCYUuF+z8/jvKmd2SzmMGqrlR/rP4Pc/oxf
deyiRc1f1ZGBBhyALmPmR5QabRf62u/2dCZ59RUx8TH8nopanEE4Z/GRKvHHVmhlXLXAMy580L4w
OlOQ7LZdLnWgJxsn27Ssf2OODD1X6uUSc2EE1Y1KVEAk8m8/lojRUZXG5qPxt85i2+S69bmCGPmB
9AXw0b2yR6J7OfyI/ZSjNInhotii3sPdOv+6m9LfcEL3nx7Ig5ODPyMpZUXbXsBJptTcgsZgBP9E
Z7a+TUH8uy/7G/K+zA7sTjelLyXqAfGWZUCqSNXkIMg4iCAsf0VM88H8zK1iu380aPuIraqQaywR
l9/qnawI/yv8cJTsYw276uUHqGJ6AbcYQ9zjIY+ovekSPbSr9rRi3dzlEXw52dEnx8auvmHX1hNW
QkemTiTtEmKReY1NJeN4EzynhOZGKWSd2cPwTnPLBp+rGkfHjIgJ9dykDPNB8UPRShaBbSctjaCw
tTdXZAgRR3Uamk6EoxBtunp0GOSOBsl/v14vCVf3EbZWlU64TWrrp1F+TzVLzc822pIE5Mr0rglm
+VOVG8uD7puzZ1DGNUcdAwIkarUZllCS9MkOgeF9Wfx+Bk9NSwDyLYvw00+YzE9FmPfHfQTina52
v/wh6eIw5T1OeBQQLmBbNwG0ohQnnqoE66T+FF5S6CvOTqGmZe7SLcKKaH+mw2+CkFLjAG6eH2xw
vtKNKffSkHHw7RdhDINogqyuYDQIAJDy0Kmz7J6jUDFLOlzifnQdmBAhGQtjuPscw+1z65PtEHfD
mJpOv7EmTlbryKWnoytZqU6WMOlmd7pUDt66PdroVt/XvFkXGoJ0FN1V9EitfP8l9hIbF1QmxDSx
px3koQdT8nHf9Oj3n4kicF6JYs3Mkn8ajju20pJ+ZF1s6XMgDPBbHrUfZAdA6hnUBUbaw0JiAoxb
4c2JOwjhQvNQEwnNrRKWPFQytj+gBEhW28Zhhe57Td6pX9qOIGUnf//UcfzpJhYDoampyrQ2qmf1
XvPA4ncEMgTEKJPuk015RfrYfRr+bSLQjpWNfQduVz09deRqm6o/I/Mcmfz2v9HaB+B3EZAp2U5j
kPH9NI3kOO7XUe0/TjaQBuTpwMijQ1D4UW7CoVh36l1/5Gq/5kPNczDusnjH/XiU75iSkyUaWbD0
urK2pFA/4S6iERjGE3Qjq6To7fpwOSQv4qzIQCFGmeVacW7mOu8YZi6cTS7+m1gBHrkm2EZctCtm
luDF9mUYazcNcc0QSHvlxoQF1321xgj8gp4cRvLNMvgPwSt0YhlWlOHXzqf67nydCs4OuyrlhIRl
ni23KYtQd/3EAWXkaVvaOiabfQ+wYPU7giu5Q2HFJmM1PfXuZ9hYXSq6gj8mgEqyjGovZ6/1N6Z2
aWN1yhegOSAo0r5H9L7NomG71GDUzFdl4WBoVCjRbSGzXuii873cQOf8L7Tn/w6bK2ljFNoRpLDf
638YCokusbv/nqJzA/DlPl4IIH68JZDjvCYcyzF/eYgk1Ly+/87juRW9VU6KwvWBNr9m5wPxF0o3
lJ91M+t/dD1JcfHGbDOcAkrYEtKqSVXzB1eGS2nkRiT17WNEtOq7zRYWLo8687yoQvKdWmXi8qVJ
R6em81Gwju9xBdM5d23TtxD1g+Zt6UxIYV4/6HjM0KIxab/MRkB9YQ+sRMaJZSpKwWMMk5nkdQGP
4/Y5yRr8dh6cp9Eh0wsvwWQwGOiA1qc4pAjRVSmNww6pJYLEMdRbfMl1b3w5a3uVxIjZjDHHaLP0
SPkwx2y5DGBPXBfizWOCLSaAKRGIbHOZgAJ4hv3gPNs7aEPW9BH9GOy2nadbGF7+1erucjGpLmON
+ZjjHfyWduczbqZH4KuI5c/l8MO38Lu4CG1HJkSDNdz9V1a4wjwYcGP/usybKK5UplU8MYPan8rT
WyEd0Aw1H8SsFmXE25ZWh5ODFOJJdVKX4n2Nb+2lx5oOAyTrLb3LEyBHsZ0EeaehsKilfUlIZK3W
Dbc1hIju4X6jf9yNGYodhBHEiNX48X97Tyc5n69Oy4cXeFwKR1isZM+MlZxxwJHPAtc86na0A8us
4RHB8en9LTsFSv+t5CZ8DkvQvGm6reMztFDH9Og0w2iGi+788wgmg6j1pF9URPtR3mPlu6olc58Y
zmHNvap+T3WIxEY2ECoDiBSEfcIXumDTPwFaVggWXVb9kYMpduTORueY42TMuPwT0MUldWlPGCTu
8quX2tpDP/5Qv4J/X3zs2QDqYZdnUNvYQFvpyNvteCmpiKtuFOaPPIkJsNIfXxgO3EKHaHoAOwmW
lu81QjFj+teEdQn8HaN1xbgqzRzFXZvzZaMw7dZ6g65b6IYQ+C9kMU4Q1fXP0Tflp/D9bfVQc65O
mjpLlbzR1JFc5kdDcfRKYrcSCLOAz40mF/Nl0IY39KReGkLv3qGTQP+3A8bH+MB/Q16PisFvKoos
MLXW6FuuwVLLN/nMUUjgAVbNFhOKp1nkHGBGwfKr7tq+mgypryF2XBo1Pmkl7JmRVaOzXo39J64G
ThxigG29+O2SZosdxSJXA7n3v0pEUBl/srql6NeRoo9siPb5eO8+Oen1rhi1S6R7aTaDBpMkj1xP
h9/M25lych4Q/bXszuRa41uweZ9VdTYPRebn+UKCi8Ly+5v2gADlPelodzCAqY76An7bSJCIdhPp
yU6DAPrRT30+qdBGDQowoZzDVM7h+8g81S6SwVSyN0A54DVfAzWF8e5IwVRGZ4YgMtgVaD/uBQqL
yKI8ZyAlFaXs826MqVHZgtkcPjoRumZBSFo07g7QAzZbq/ES1CjE1KErwmBVir/mcmpyZoxLAPGp
uRdQ8oveiNCEhKh7rfpNISOqksEVhe3ygXXg9AhYyvh/rtnp9IFrJevyL2pgWomvmQASf0gic5bQ
6xnBTxx70XUBRRd47hzggdMdbZaFvqisuQZkAMQl2sAFWc6m5Zem5y+bybnnY/wgj5MENHN1KTlr
Tvl77RdV6r+ceRku2WvS3aaL1BxevCFlS8Hb5AmWDyKYduZGjyHU9oxgVebueZxWqYatwSc6TprA
xab79doGyBQgBbgsNSTsyrqL9zRprDQ9XcSGYJqfz9ibam0HayF3vQC2evPvYGsaNDXAH2qAuzSs
YBYaaXBtqQ9Tw1QohjKt9MbGWE3oCdRUgu8qjsRiaTm+vIDLXU93cfCNY3jyGMhNACkjiJTrYeQv
NOpppvF+gUxLSm05nULMVwF79q5gB5ZpV/8Vj31sVzknql8NgF7JzE8ab77JC3oZoy2F1bPT4lwc
HY6qrs2kPqHkfhRwVTsKVVObKPs7Sh+LbkudustpTghSW5D1SFIqr5cfZC3vVbcgbu/wHphEOtQX
Q6WfVJbKidJ8uvqBmsc1r1vLnO958ccZv9PlhU7/J8B9TZ0rhjVJ+m1OT/4M55ew8OjqEXO1QJO1
5BcqfOmKi7Widbcvsrb4HT4kRvWq6BlWXu9ELXDoPkHINxoQxdC64C+xAoAErboqiGKPDDxHIhe2
183lltUJwiEB/p3ozHmOsajyYKxygujRgfcomJMKMwEe1AiEPI5CTwP9OepX1GdYJrqLeVs/QzYo
5rsNcVS+4j6Ois9nz5AZaS/tl7wFc4VleLk2bT6lkZ6sqXMwu3VN9+NSgiKmkPMdIO21YwaKImfR
BDTnMTlOefnONF/bKnAya5yG/SWMI0YqyrdrNNOMyalCKodaOY0RqZQ6xuqvdmDpmzVsy8mkOnyZ
JBSGkU+kS8POmlcnhSzYPxr0vPy6LhNe00P5tO2H0cnRX82GcAG3UxZVuXK1yk3vZ7UHGFUON208
w6VxdySQpJNYSn2FU3q30+Y3T8PnKMnj7hBUNjnaibzi78Pns9QQ8nSfgxt+AJ5G6ZBFDCAdR4Ch
3siWToOcujD1L44BRJnjj0m9usWfJT0dW6S/gexVkEIGTaB8HMN+qvXPWh5COmNPzEAPIxVNywDn
T402mtXw1C0Y7DiYVPrKIaTSi93qTYAKNUQhZhizVYFWuk4PzoPHFUHvgjSaesQkU31TruDLNIUV
qvshZvWyDDyYqsOneKBEsxas+CmopPVDw5yiGokHL/j0VAQZCQhSndxrHgE1f5RpVRFa6tcr45e9
+eg+Y62qk303iMLqt2PzSg5kNBJzY4I6yVsdKqkPL+PS+HTt/nfFFTZL6PCavYt4qZdbRoDwnZeq
o+az9Lke5sOgOc6fB5i2ZpBENLbHl5O1efpetIG+cJwSh51OifTTXsSDrQilrGjEbiquwHf03r9n
Xl63Kx+Wpeujb3AjHCVOJSE12UqQrBc566BHjnoAxKMxGyMywmrE1spG8UJ+/8mMtaVfF1KeRxJM
vwtl71SD6k8MWmCrLxHDKCm73HHe3GJE8TW7XiPggaDCXyyt9wDGSenU84eXWuciGm7cL52x8Fco
TEtSpOVxWABSDLcOj6ad/lbHv8FvAA4PAylhBsGdcyO+IJbs+VWtkaU8TY3hdYYFsO0LF6WgLEnL
B006bmX68xX1weXZgNwGedA3p+OfcsbIPn3jEnPmHFCsnHZddpkxq5hTsZSmdUck3ywyPJz22Jp7
rF2156Em/yOYCg7J6uXj/oESKzYNrOngUiWiH+f04x8G+LYGi1jePzNw5bpH0iIq2f84PwsaG3zw
4kjwI1tvGm22HhfWNFITNWGhmEWZPZnVh3GgSr/xaIzCNy7dzko5fbQ6696NbeHzLy4iFzL0AORt
rd/zOKhvi/BEHsA3lxwRVfc8oq8F+YiXIGLN+x0KmQMEemJfR0Xb6C7efSisdDBQQ4+PCNfBz1yy
FrPgu+XQJfDPYAyZc3ywyl5vsIcIQbRZWBPLpxsbRK/CkBAqk7JMHLiByGit2TShXLy9YmNwXotc
7KkMQTP84z2mdX6a23EljVIj1aGqUNHgfrbTGTHnuteEcxNjvhbukTTzdpUFrzWGstcka7PTZuQx
9lk1cCkENv4EwSDKCBvG4wwisuIF6XHkA/qtfOlBHGjpuV0HvV9hUZ+EYj5pXSkjRkckk+Y2fVpI
hrBr/csP6TiWNG/J7CjF9g8SiCs0X8xsseUawNmLaqj/7+8pehnulGjB4vCeiOdEnAdINbBvHHZA
Lt784TQVLa9l9c/+pG0m75qKrd+VRCOPYqy0LpIktPPBtLhatt7k7D0EkU1YPj817TkBPyMifKlJ
KAMlq49Pb3P7+vf4/WOm75z7GvXF7OE2DypBCjEVux+cIaPWEq8Fg+krHddUT1DX4nywU+I6/976
0zN0y7VwOnqbjKap/foZhvj+TsRcOixGSwlndceyMmq51iKnjEuzq9N9+Y7BmoHGohdvypIHhtAS
sIogrDkmm1fBdn1VG488/0o6e5TGdf6xX6zyL0VhDOMFAAoRfl8yBZkKQRzkv46CKJWLawTeykUl
5HJ/GTzRlsT/JVxLq3I7hFotM8erESrW+PhZDbXWveIqwwYnDYr3qbyj8y+/OFBH5w/ghFsdF4pR
jwfA3VW1vC4JAK5HhSR/dVpWRq7B3Q9sF9qEdrvY2ODZ3vnAruRas+msbwfxwfj9KD7kksbmpmmB
X9si1UpVfsBEJmbk06nlLi0Xc2hcQteZsuYKi6OdWfw/OIZ6XNtdzcsXd8Y9svPL/w7gIMw/k714
doom4JfHP5pnRLqqh/uX7VVt5mSIsJCN8qwQtRwn1NmNEA0hlLKVIMlJpVtenMJ4u7+c6WEXcUnb
81avZO2Ub2+CYmKML+JqoCd6yEIASa+yLF+30gLF+neFBumHfcBi5dYfs550oWIDseJUe/qMy+h1
t4cqH//93AToFcWmezprR7VZFwGz/j2GPBfV1B/4tpMmrOxg/O9hhZPKpDONArSj4NDjeg6T6BCE
R53lwLZuURQHws/VsC3wl1EcmWvzt3tQI5NUk6079ThNDvxS/5IcvragbSh5Mcs5SLCydUH7GTig
YOU8H63iQSawwGfx+okY09/hkiahVcAuqei2RnvGtJb7iyD0RgHnVYdpewT1sBFpGHEZJAPImgSC
TNMv2FFCTOeUaDztNPr0rLZvtY8usSIGE/97Nn3Lm0UEabrVMsZrWEoSiRnY18+R2MFPPad2Kxfu
Bv83FpL1jCuUPHjZEbRENWbtJH1OFAlYkxMl8yRUti29yTWg2iNYqk+oE3LpcMsRabbehURWbvdx
5YVkurU5U6h0bk0+p2llVdWrG46mFSzspTcbuECE6P1km0Locc9aE7hUb5wHEm3moVyhNfAuBpMB
8PYT0YMvLcG4VZ2xlap4r3qOjQ4hUReD7mx75jsOEyACsVNKKpER0XEbb4xyfr85uNJfnz2Vxdzq
97hbTEMsc12ZolGWQwVXTpPdUNhQ2SlK9ayZLmzIPvoNluOOEkSzOE29Orra4L+9eHBFudg62pdU
KVA79SJ7nai+p5Nl/ZW7qfFPq6Nw+Oij3vOgCZJ1x/qHjnzf3h89Faxu0CJuUjK53CHS7BBpXLKH
k8YWmvD7gd7LudfyFKMlD1g4VlG/QiLaokCg4yV/lyF3LPmnUIMMl0GhZ57jw9j5NNSXyr6eagX9
ksdAktNAkNu6XfwOmU/4G56HRiHBUshTfFY7o5JSDYjsZKkm4ofGbq0dR+L9OTBTmGUS/RosqAbP
4myilLcqqzlAcfJMFsSIn329ybPsKP9PjcEuu/LUhL9Ug8nn64OIwM1cRulFXDPfkJOj2N76CV/z
YIv3WcUbw5PVuYyZAN3ozkONnDpXNAprL3q2qV4mZDLEI1ux7tl2ftT6aydtUXV7K37BWs/95he/
dyMEteOhQNz+JeGZi30/dEdoIWf3vbjN4L/kbSTFL9ZxPTJZk2NjH8m0ieSEE3LDEYXlI2q3c28O
snj07hTpqHnQaQK5f1SjsqL6cH+wSJytDxUR4A1Q4/qM/S/10THaaI81MA4YukPyLQEZho8jIAMi
nBKkAxJQDoMCDie0p7CbEuhyKEjSw/gC148h93pI6ISKKVkj1r1POjSJeIzvKqLMOd7jtqDUgU69
LSDMR1/Uv8Y1KSMxxJMO/38eOnkLBusCs5D8JDSRco2XYoW8dp9pfDO1ck/LgnD6KbldU1u2TkxU
RVgYMXQsMU4CuYVwQOJwpnH3dNlLZxnV7M69IDP+iw23kSY9m/oDH+J9hpMfLbsfcS7TbFVR4sTa
UGRrqzPbl+/VZasimq7QMNcGlftfNS3ZZRAAzIFrlUebe43DDCrnGPyYD3wA1IQxVdSdiYaOf3zr
JTowNRHaPZLNUESjdF7ZFV/HiFyAEjH6o+uOaaRZrq4EbyXe4gEj0ee8dwfcfRNvu5+1/Iy5DXiN
ZLWAfRAyzdp71Q3uoJfw2ajo4ZAVvwEarIBsGpkGL+LIdYeBEF9kJnxKK7TkY8RxfSz12w8P1+XB
33y3Fa92eGc1UnXZCt+upchxeu9ZpGCVoO+3AzhiLtQ2T9jrizEDacu6SUx0yNgXO2OqzrCkoO02
wAwGSMVxbVPBfKj7psx2zEP0xoSYls7i3APp+nmEyqBBytUghzWBoKXo07y0QjETk7xcLetX71MT
sZLKm2WUqRLbHmw26lEr6c1TADIVMBRxQ0hUNQyMIfvVhlpujVj3Ag4ht/bshMnzeinBo4oJU337
GZMlQH5pVIJ7wzx5wI6zgeUdTRTH6PVKG87jdoXQUusUBigTZFWQIguPlMydTHajhCiN8Dnlso3e
zKK5HENuKUjd+ZyRfQ2lmjNEGVurc6j8u1KAg1/N3BkSqU0FEJwTHdGrlvjHiR3Zb2LhZvNRq8zU
X92JCVga/Hun1uJsAdXP2naqDKTursN05Y6JZcNP+UGIcSPmxQU5pC4oUyDqwF4tkJJm8TWo7wHY
hxrCAVMDZMFYSQ6NapPLdte/vZPfm0tnK/3EnREa6GzVM4WryX+YnI0T12py5PafI3rEg6tHxSS2
0CwZ8M/pbOw6YMxbZqYB2pVw/JFfTsYrTGUe0MFFmzdbgNVf4laWQvSv9fu77sfeA5XzdWveKbuf
m4C6iDLU2s2jx2942vMi5Pd1JkqRrJ+m2ZjqWfMErF1FavIv4YFP9v1wJVX8r9yShOL/kUF4xZSW
f0FaqtbiKMFXDba9ETZwup1wZO7Q4RtWBPwl2X9imxgt9jxy1o3LgpEbI7ogzoSaQlsNj2a6NpnA
q/qTsyJZBlLYBFKhNPhVPDNTu1SYhQ6G0ZO4VjbZUYxxlsmiuAMum4lbTkReZaJR6ysY9yJftGKf
Syczw89jEcl35wwk1WP/rPfihaCTlW0rFWbeIvWzJNeTeSw7wvacObwNIldgVI4R0xU5EUOyT50U
Xfr7NXuCr9EVwLVkHewNKPx7IxkXqCKzgpFN7BLesQFUmgfgES9ne4dmBlEl6OB8gCISFXDPpYWb
gK5PW+BMmrrptWFbpNqjsPZOcIrknTrtqdAD8skY7539XmTQwci9fndQKsJqlVNMedV6Ljb0Gqle
zHnAF3vW+QYuH3iDLvK463TswFEzOOBgCIDMr7/96FYzOvuHP5EtTJPGK0vAGwgeNTj/QYTW0Nkv
2F2Y7qEnTYwVb/Ju+qgdazqj6OCToeH6ZnzIRiirPBDjaBi5IKry6pYjOZRwtjg5Vb6xI5+KGHFc
OHS39zpgO7Zg3dhXatWA8hsTnUdyD7SgSiul60tB/hSjJq0cTU/UQcDdmGD3+mY5054myLcfhphc
KdUfp3q4HR8eBYBBjiFt0o4FY5mnMTctIdYcbAhKZ49MN2arUokbSCKbXp8Zsey8LbKb782LuULz
32FTnqwnJI9tXcCBR3OfzM0jdz1YLvUrMlf/wI+ICD9gXrxTdKptRkj5tk6r1CHFF/XcrUuOpOZ8
jlLCDj10SvJhXCBROqF50qQaXz4X46YRkNljCdPFLQr/SynIxrs+JYNLMMiuv39d6w60BBk91MJ3
Foyohw8TuYBdMNnz34wwqUfqvMJVhlN+LBN2fnvdKJ5GDqLMDBmSDCDAQ309nfsOvAGFt0/5kkeO
cdKhIAA9p9HTx2vOkeb9mRwV4LU8ESVCtJ65AGUXrDdkmExpw+VHQpgRi4+NU5CUZAkVoNtsGi+Q
I53JKsmrGXdksXE2yJbn3ZLUAo8i4Dg8hobkGGN8VYhm+XkJ8BfHVwWEreVCYH+sOVF5NzJLr4F5
JipIJpLSfGJYfaooZtwsNWn/lNhIMxklXWk4Ha9LE1ZXfqNco2MqIv0lg2kH5J822biEa8vYAyYu
jnprUGn4gDtGW9HmEFnYHMllqbv0bQEttxTJ/EaTePGqI5Dz3X1j2ay+LiDrmrfkfcsO7Mw18uRn
7wjiyV6ohcbbuQ/bOP5AmdPt6qvsgfAiCn3aSnDnawRgHu8vbia2zkMms1/SElhC2csYpBi365ER
DZrK3zED3xY+3VlhyWeQfh0NrKJEe2a2lKRfrI2Ijr8a/s688S8Pfi1EWM+MuCl7tNDrQdg1rlMH
kdi8NslJSDzP/08FPh6lQhDQnXUNmCr3bz07D7kOp/eSTwMw96hTM6fb7PO6xC5JaDHMSB6XTe70
mct6SUJL8z9WJNaqe+5Kodscs7k8/IPKDj4IlH/UC4mFnkQQeT80imwsQV3H2Gic3LRKoyc0HG4D
/dOzxXF+fF1VNhc8FUBE5F1uhAClDWiSgj4pP7jvlnrm18rbBDfED/jFgQVKTrlDbWcy8FDy39+o
ALkv8FqkGP4+rc1WyRQCLfzuxwlCoCI9Bcc12YrIKERPhtEPtkuT1JQlcEkFZTvcK8YZ/YazJUNW
DShJYAOXMZieR0MNTcr2KBNYmaPNn9norhTbLTqQPLln6lldTuAtKmDiem6siEK+taqljR17BYGy
wCpTZCcfr2DvEia4chQAp73lzXySe8M4D30nJ25nyfN44kjsLcIltJ3afmgja7jXIHiNSztCYJe8
oFcyPt6pv1mrbeNKDEfJYYhVP6nqKqr+h9yfiQ/H5INL0PcvprpGj29ydoJ0ugxa7I9vbTk2mjEY
DS+FC/gFQAsJroCuPQB+gFgUPT9L0YCyPpA576aaUPYarWArOyPXg4xRVMwhI7p6lpXXBbb9fDxc
iALNDJnmKJbavFukkE53U2/483GqPrFxnHnD2xRut2VxUKgdS+//aRHdSPRLJr7+o0DUGW0QzJqc
f2SVt7YU8or6qXH9hdIFAQin9jKwJ2HSaVikhwHxjUg8JfXL3nEBc5rFVBhIB3HaaoLQg6kb9E6v
qdcGVyJ4qBVsFbVooJs8efDrLZ92q+bEL4nVFfDAoQbWXW0c24m2zHh4FF+sKhdWw5CcSmFDZ9KC
7FwDF88dUK9q76vV0e3Mvo/CrYGiT4Al4MppJKoPK6Dk3WLhGbVLgbfCF/3GQ6uH1LP0UNRQdN3z
mg4vodTUMCUFb7IP0ROAv4BS/hBneN/ZyjR0byCery3tXm12yCqLUQSmvTBMLTppToRe1mZ2uIxJ
ApXYh+xL2Bxge0hmUw526aE0ImisXR5KOjL1WJo1OJN6QcS+QEkheQ+iI3SdAANajDTeQpkuptGI
N0Nz/EtP4jC06+3k7IGIG1F5vTGXX2+7xKr7C5q2gjp1xp4pDRO7kVHcQ1oF9A2W/ztYYSeb9l0f
sINBW93wS8qZ5ismfHej4+cF99Iir9OoDWoH4OwPfwelpk6vCl5KU+F9XCjo47xBvoyXQ09//AK1
duc9C/6R8294l4hqCL1DlukR/s1qlHs1Y1jqNatSJYC5przgxo977aGD4KXGHx6cdGT2NZv9sAFf
G2AEFM2P6ObkpOf+ERo/tBqYtv+Z+GPnlzESQjaFl2UyaAWVMlGStpgiCBav9JTWwGfGdz2bqp8o
5ij6NgRAkBU7Wbtlzzoez13ZAx+ICqKh648O0IywkytuIb+xIZwcACe0wHHZl5QUnj44QJoWu4VY
3272KewiVXJbLUN2eq9eI3H61EAsj7AvXNbyiEuxzzFAMTW4dgk79pCrgjyerQpVt9yyXJfvDPDL
MbSi1k1LyDNiScpMC3rZ1r33xGmtbCN/X4AO/NRKz/7/SbamalTy8oFa3Es0UE+RYPtuYzwuBZFQ
6i/DVAStHv7LHdyy7AmjZ0Tb1XSrKXU4weXxaJg29lNXTBNecmWsmMlh/LpcD00HKpwQFMtqpnyc
j3Ie4SAy84ysmveNaiqqc45lqGeYS07Q80RnlHlfWZbTzh+SfJ7ETKH8twHh7q/od0x4kGhMF953
zM2SgHVnbLlR2cAYK32ifprUgRalqSmNUxNdPs2ULzKhSj35mQz2FLzG5T81pkWhtsgfaVdC70c9
1b/FmSuaLHpPsWSjW3h351Qb0DJxr2zy1uftZj9m4T/Dx+iO8yCTOSvQJrqsvvukfoN7euDuv2Rn
AzmZ9wxsHAtvLTGN5LtH1q2Ryt3NLK1s+P7wdd3XQV8PQ3qeeyv26kt9PKd/P3wGPTaz3adn9Qaa
+jNdMS1oI8YXHI9ewskopjbUSYEzwA4H6A37VAcLSJmr+OD22Hz2Tq8upQDSF5BIRF7+3DLFMYrH
RDnIZRSYxPl3gpYeImLTiTte5cJ1xooq464GaKQB576BKUrD9JgyP8dySdOCzVpJ+KFK2uxVOLUT
Q5r5ZJvUn3M9ODWIudoJDjGcPGJ3tftDIwLHbYK04QW6KoLLEEFTpgdLk68bHUjW1o16DNl/wFPn
8X5YwdRoVPEvL/4mcoqEhToj8yhVrj6OAR3/OYswanRbX3DXAvhdPDikZXT5JUpJuIq9iSowI54C
sHw8xskRPsvNk5i/4iFurC0UygGgHbjeS3OI3D6QSXRDQzZCLApVU5qLiMux8n9/p/0zZi3HGtRo
deZph+yg+McEf9xeshm5e9k0EhnBsS2r76yScamwBNhSvPHNdp9EDqTtUDa3oIrzDX2HqUL5OwrN
Gp9ju2qzEPwy4OHnv9VXSj8SJSJQosM7WE4mho9VkVqbZFlXvYDZqC6mYcLWZjQjf8jDAjkNOE7E
uA4viDMUl7by0twLbdiXLzjEXjxjl1L3It4o8Z1F4gvhG9mQ4ypy3tBdg+0t6v0/+c1oBp6DgtKa
KJOpdytyUfT8edypcDidh7rtKMaCL6AJKQoF9Ai1ZldokNxzLl0vNUETTUFZCCUXzBhTcJziu+Vf
ZkzA2Rj7eOI0xd6QPc5t8O4YHxV55qMdaBNufJwOT0a351nccSYxqgOpJPd9Ge8QlI+rYtz0lD02
ijd0rjDchsS8q5dbSiZKKHHcT/LmM9frN9sv7o9jJPVKCLxLDI/yzRnm40Bw9IK3H9oF+sY6/KWa
ABQxsQJK6RGci4IikuXJa/4tzcNBjIZ8f0zmKPikJclvsDoDHaBaACKIrXqFlTOTw/9o9aguDsJm
NR0E2oToCAwY8pVpL9uQ+F0E0geSjf5mXamTbXa1SJx2Up2p49640dg4i1hOSlzhv0tTF5y1u7Zm
RAW4N7nFmwmt3/iKllBTehsBgthBlqddb7Es5I5Ue4D3weiEQYx5CFRQUdSXjS5eqcMac/bpoz35
hFwCe1dsVRxNMpyic5DfV9kla/dmBgBaF5Kv70WNC/Rmp3QuUtp3o6H0QlydWdjGpJVSzJ/8BLX6
jIAUQKgkHPZoRZCN+/IQaBBqF4MtJqRIPeC/5wfG1Ud3FYxt8CK8Sq6X1B6086zd0J6OMK4KtiNU
fH4ZLIvQSEWVZEbyzYSwYlTzgZZ1oW2/wKrimJwmgJrR+oqBfyF8HRgdortiH2UF+BjKb2wz4fmN
enr5ActP6FUjLEIHgOcMY9uWaZWVYvX3gkXurwx/YX5MmEgntva+eByUNbMAkoccYYXnFd3YawNj
Y8j5Nnj8D5xLTJeV88mrmCVaRp/QIf0WJjkeQfIevdX+eKnnsxnyuDWblnhuwRWFpQSIXHJarfMQ
I6vvrtPJTlJVFYt5Nq2Q+wmR1mCzngeL8OnMsV1oNQyHlMAuWJel5ZJin5Kj3uJQfgthmhVEQWfS
F5H9Z7T6xjgk7NZW/y4gbiaX3wmqq9oZ4E/nG+IlaacUxuG8nETsSxM+zj269H5MwoaQudiE+Gpi
5WfU901uDifpZg8C/uxukU7tg5kvduY8tT4AjC6/UxXacU0w4vYFzBmyxWizxZTN7zC5gBD2BaVx
MhZtyibZGlqrlpTy93lvXJ967LGmZU1SVOqDIkK1I36FuNzIYiAIcB1xHg4AVP34w2vM3Vr52xEL
L4KW9KbITMVb7FTEhTI8A9BhWYka8fQVHagmqAyJFmtsSNBazpxBCMSVHNE305pXAf4DoGd0AJoS
cs7WxeI3PmnBqqncs9U6ejD+OpdjlyWnN2VFwf+rlloyFc6U9JJBpmcVchgzi1f1QmbzirJpex8I
QYR4zpIsclnot+g5xV73dCEZetO6PSJh45TUFQpKZrscX3oSJPraS68Poh1zCovE5YqBUbSUNQJS
ptTSa1y62cMuuiY1s6UQljki0ZlVrM/xi7QVK4lMETa+ZphfH1obF2d7QuYK34T1R38zQMIzZpt+
UpUrzBAUPVDg/MQtxELeog4sOJLgRUpZ8eaoGcwnSd5zAsZOA2SjBd3Oq6vyVXKmSbxssPxSbPBQ
qE8iXyL/czOfm91BXzNitLVIZOObQJ/QoKZ3+oONi6LiKV1qCRBQiYpI3CTxTp5OUCaMoWdCnNc8
/Z98hHMQD773bAe0woOFteO1NDIaWM8Jqcwg/9jhoU5soIOVifHujM+QXWDNTMRrheKvSAm+TnoZ
yfchgRKpPYWaAH1uA6tFJCdE7PeyjgAsfAr27zwhP+Tf//UXkzxF55YFbsl+sbHkcdjKJHjBIGHl
I6zK5/8DijM/6dFTcb4D4jbfqGQ0GMgk20BvjbKBvZRsSWr8+mQ36cKXr7v0h/3qB2Iuq6UVxjHe
Kkhhpy3ID0rs5xFNHWaELsXdzphnAQiVGLKL+OANO3HxWWDPD5bsRbvjsxDPDIlEuZ5GVarYXR4p
rgNoa6l4AXggiUutm8pw7YtFij8uy94P56K8chGEn+J8iEqT7JRxcdmDCNz7xb5htdplOSup4rUA
zgMw0awUikzdRSL63XCTwPF40GmSOExAekORTjp1hAyYdAvPxjBtv+H4+PfQ+AedOtIHf1IPvKAP
wYMLRQgz+MCAr3J1uVkv15NYCisQAwsAWIDg5NoI4c135ayRhRcLank+vn47J5LSeD6z3pZ0ThsY
KBCagqmpWoo/X2MxcmaZ5ub4vVDLfwNg2EbwiNCr9TFlWXdMzS+5O5xM/0giAIBKoU8Q18U01jg1
DXXjCXYP2hnXcxycNkfYajQu5YPnSpt+W9ezmlC9YoGlLZ/34XW1QcnMQ+oGCs+Y8WxH7wtwvrj+
lyOGbF/0Vhpriz7IKlFeGFmyMRlNjsVuOs8pVHNekuqsNgtjK5GEzNPncQ4lMhghgPR4wJ7054mR
I7Sp3VqP3joEYxIQS8hOQOZyQwSQ1fLCsKGOoACE9b0/zpqouoLBeH6bif7rz2gxEHq0SAbDueJq
/pUnIoV2msQC9F4rPkwXHGQwpmJiPAFGwj5vlP0UvRpPbdQROysz7TXTfL/c2xuZdrqwSMHk4kUW
XGBHu8qqyrBKEgeffpKynfKd8zTV7Uu+Lnri4PR4ivyXO7cs9qeV744GNc0ItsZ+X4zxM1UTUy6M
wSH3naOcNWSpZeN8HXIC9YwLx1o4QGq1PYvCtphPiwFAKnLtIX+PPHHBi9GhhPjZbSWhp0C9Zbjx
CsA3k6L7uDxaIbER3pdHfwUjxQHmB4NFlzBp8j5wc+S7H2xhgVTTEK4kJsvF+JGCbubm/mk0oBNc
sNPSu4fNFU75Dn6O9EeioqJyfOSapdsFNEbVpHUuUpNQHBaBzUscY9mCHguV8RtS0WlXXiOyiB5Y
Z/3HPYpuHVwcXN2qpgF8SrX/EOxSx3iFGthTxC48XLQ5xSBp4XhgmiZgZNod9bdxXlVvLCo+rkS9
MOqXHwr36Bd4/8Gl/jnD3AwBkDFBBjblInMKpIWHWmeBXWBLTQbsowmV2HbVlM7V90LvSy1mFKiX
9OklMdsG2dZWYdl4SIrUFrq6GtIPNLdYhpM4qiY3tfnFDIM9UANVea2bS5bo//MsUSv0l2y/gEa4
bayYROZQA+ojfV2gsHf/8aBbnUz+bcZbUrTODjKfrKI/tBANOe3ITb/QzhGDt0r+ktLOpWvoanYf
UuZGg5/GM2TCQLNufkH05VFa1MZJb8wubWN/maVmMmdSmZnplfrmj2GKwOJ+YdsUTXoOo/Q2l/Tv
magCVy48bcuH7+AvkNG8pFmoywxKJDPA4aYld/QXeijCnV5fgB22hk0+urOYm/W+5QW/aZztAHq2
apDhn8IpaBkmjU+XsSOolj1pbx2COtOq7mgu7PFJCZYY0U7kwHLHNUM812Gu+JxdJm/DjRvVueiu
EfGI+aIpXGLy1HPPNiLv92uwBq47TJPx/IIOs7fu0rYD7szdrC3K/4UPvwqqkysNjZ3ciFUp5qOy
y/v52EEXGFYpbgIFn05Qb/RpWGb/Un7ccZlWEqQFV4QZOuqvvlxIBFx3dX1YuWc2ChZuy7QTAz66
p6aDYLUjljaOyK8H7oFFfPXKcgNJyadxPzI/ksQX/rbuL//oyk4G0Y2ig7qxYo99+SYeYGVYly1B
0OtgqCIxrQWgks6o3VqA2ejvojt7kSUlxOq17l7t9z8JYp6Mzapij8dZy4TAkxFr+bkGymJ6+/bp
4U//hD0Tie46nGos1/GhYDrczbFEdImuSUZHPXJaG174vZRMdJsoUXFLJw6ck2uOo5Du24BHYo0s
9WTWrwB1jiizA2g1wo7ONSAT0O/JJQ43rvgNLzbEUmKGsryZQ6EQvCaMxUuLNX3M+ms1vmJ+BTJJ
bPuFMsmKwA6GQaPxNWr0mKBfB7XHo4wx+L1ER2qn1yJUww/augt+FxRFjGnjgudQbExKjYBhMr4x
q5i2RCUod5CNNsY8YuDl4BmAutwaPgoUirUKKIUAWQmHDi9Qkw7KNYOrfTrFY584UVNDRhyBZjHq
ZDoa5W2oT4MdQDsfmtliKd7+C5giLNRUrTvzeXM5LSMJBFUGrIZ7XvsID9hdNcBCnKISID5HTr/d
9Zrs5pYC2q1VJlgfKUMxvwKkYUjqojPSgPsaBbNZpZZX+yZz3VCijbQWPeFSb61PCrdzasIMHTnk
9TxLq+8Bif5dL3nPmyBkbv9f0dqOhkHr93xVQel2LEtmYPIqFya81HeP6f148cBfqPa+V+WHCY0R
EQV3O6J7AlAp2CJaTSdUU47nqvQLqh/oc/KrBCDFcLWqqZUE+e69nzA+CGYohIyb8Quk5oZ2BYg0
mIuDxihNJlnBjLE4BgEGGcFX+7g+EVxhiFnOmMo20zPOMzz9XR6TIbnJJ/ngIIL2rJoMFs6rax+Z
3MOWNVlwuArsHjths/AVl9Ff7bEPxqwhmPHhYNrXAW3/eYiVXgPhC7FZaP8rLDJ57Yh20MGLina2
2XLbxAkMtjLvLr1+konM0bfwQgJNtF9M2UwJDYU8lZjTNyIFKVYWvUSET8GCnmpzeJxenrtSk/QU
c08gtrvX2Hov0ATcHgkIzEIGrmmajZ1lMOH+P2/iVEe3QVdv22JCilDijiv76mdF2x19cN6m8Nap
MPs6v52ORpOwFgTrPMIdIO9HsijVh4t111Q12EUkVSC2l+4UetcRfxn5QbQXkCp0GyCjxtmRwUfO
piuLCIYBSpUCpSzJg4tOS3HQDJvwJbeleRucKgWMMvYkYgWkxOnBZarnGTrPkodGbC91cgvmir6g
KtEhDVgKLFfnZUEU7BjcYkkB4w29bq7XwM0GRWxyftDkE4PvrmxNo10LkIHl02YKePfFs4XH3Vz+
8kymz97JNWzKbtXnUAH34I+MzGZMkF77OYYgb613bHWdQ6wGh2oBSn8x7lL7Qgga06a9BNoK66xw
3wJyuIx2N5+5776F+TJjZyTHyIM5fmncfmPP4SzmvGG7F+KFDIhfhnZrrNkBl/VHOyoCrNtUKxaC
sibU/4tRg3+RRo5qZKc0rXxBqOGnS6VCLrhZT0A3eQeFrBpTOzFKbIRJD4XDwjCrcwYzuO85Pga0
7VxvdV9+RGNX9rsKM84SGHExY5sW+xG7SsLeyhRrBxAPk73Stzupd5DbxQ3fZpFsILw4btN3/J0Z
fbSkbkT6AKCTSg/KlI1q9FftOCgb3Mdb1U+2cYd8LEOQ0e/VCZzfxYK5Rty8+lQrY7kfK48f/Aod
Rskxn0VSXyO38gRnCpOYD1sA7n85GsZGIHd3db5vNO0d3dq8TbiYZR/Ezmf40HJHa3ohkNaPn12d
6eyZNRrZSrO28vtbqo9P2A2yy1zIi4BR5nfU2MtoTPp8XFAxssKfmUhBg+U78e/SlM7CH3AQvF4D
ula+oVuLrl9VXt38KP1m0JadSnYZsg1H7FUTITouXxwQ1NWQWh1TdTuKcXxj3lyMffG+QKb6omFp
wFsmx18qMW0nPjXO8i7jnDPgT3yhkioaTrZlaxWLYBkPG6sddop+AF6dJQU8uVzUw4x/hFSaPKAT
Sgk95nWShdYw+Lojpdu6AULk2m7Db7CnrK2QEaOoTzP6JxP83yfGRJOmBqJQzL+8Q4a1D+5xRHaW
3Ee/aJ3FTb2yeDqmFvy2kLj+Qap3S/TwHMsUlAtq1eHGzA/cC7bG3+PrpOcTEXC51wOnZp9tPJyy
T+mnfsISdnxWYJ/UNuFGJw3gVydhX1VBwCUx5wxYdNgrU1OLkEhNor5Pt/MuxDkyU1Ukq/AVzmBi
Zq6ymbdG6bxSUCBDLHTI3D/gSWgPshCBZPE48/w7KBIpE1iffKa3qNvcsM4rm+TRxvGooVmSnoXT
sMUHY77VqI2UeZuYi3ha81eLTB7HwwvVbBH3FGwfehtcZ6Ds5BRrBmUACpdyHJB64xQZYSegq0oB
gTIjd98xKTanU4kTFphrnZ7n9ufzn8xTc/RvwcPKcFU31P5+PykJTQpjWO5wTD2FTXPAWuRd49OZ
F3WyQP+BWa1KosXcwKzCLonC7D0QLEoulhh4vlFeVfBF7MAyYDCDgnTeXuur8NyECBbwBn31EBB1
kGIqRh7ISU5Bt9n4CWmGD0DJUPGXTqvHi8y3NqINtUu1Vh2Ob+aZ/AdUV3jkojdeYf6rXVJst3tq
/cVYIx0IoUlIbUBWazK+0XTTnOouA22wdUI0GPjXudUP3SRzQxiqy4sNgVQvWMIgvHaKjDYVoHo/
qaRPccAt7ChGQIj8vYn2e3nCU2CtCuibcFMIRYEqihdtNMeTxZN061bRrZPpYJDilXSYQzZJz4Ba
Iujnj3a9boL0KkysG2VzMBuz0z3uZsCgicyu8IF8FeBNMeulQi+IaJcTKvyT597wvr9ioCliMEbe
bMEB9NJFG8ght0baaaeVKFkp82bTI2y/HinYEBxoGKsgtBmJx0aRoFlgbg3TjXL5cF+s6XUrIU6C
seyoOt9yPgbrdQ4Y47qOPUQohL0bIZ1uccLGcRye4wbCFB8XsI+3z+OdizC2jVGG5mCXBihSFjYz
slEzpE6zzck3qX503ADgOc6hrL6AFVpR/gk/kDMBwucfFO2oNWAUH+5e1K/o9g4r/8+KcdzGEfjJ
ZVPOPUCNApo39bT3jDZ/ScxsqdFz+a9Z3iT5VFM56VDwmFt13DRuBLkBVVB/6qENIlz7o1Egucw5
w2RKh+1h9FyyaR2U34F9EXBrFQshMomkbz2CdLybGy7Zb423np6yHZHfxjnbOrw0foJ4XMJMsAee
HAsDDbimO1DszdZHs7CjNBGOqRaeHaeiYtiFIaSzvPlQU6YsZbadxwl1aJQVZ2K4UR/OUbNyDOH5
dUyGqafMQ7BJyPEqF/nYDC8PMUNvcxhebRniqnb3D+cXwwQ4hU2l0dug7pAfWdrV0SBmTSas/l5g
e9Z9ZD21OFrFnSNx5W5nDGqDmFGUte198co7ahZkQ+/hCTvIJEy/AKz279A2ZInUhraCMhaTnRmR
l25BbsEUsHt95vDhPFUH8HvL4jRfRTd2SCQYzyTkGnvyS3DPQwvkdljakOWPUebUozoZn46qQKZm
rRZefX6Y1Z1n/HCG8KYypkGg+6SQrCAW1Iflk/9lqwvkkee3XsDIr0Ee936X5J4KibLSfSHyEC+a
UoCO3YONuiS/VyKzZBv0OZWC8i/yJTXvibOWpTZzEg/DzOQNFf6mUfitHhH4fv4JpjjJCmUgbkQx
XR7v6fxSSsYJlOxlEl05nFzw48BrTV8yE1NfNpqbCduKZ5SR1deP269GDbaCx1SeQVIJAOxJFX83
3M2JUsV823lNWJCMm6lQ9w5cgkOuOjlFCpIE2+GxddjBZ0rkqTAJqMb4D3RDZFLF5PQajO/FLlou
9RyJHZkMzBT40o3tq/h0mZJiqVVWUU7IAXYqK8o1AwtfgE2vhqNyqmB18myNctLLny2bi7nkjOOU
MYSyfemUFCeDh/l4ySO7fBIGR5xPxYjrgwhjkZKYQQT0HiEycpQ2WXLVveu3ExAznbnMMF8AgbxY
qS1BQ5BSq7IQrl8EXGgGTVdmTWSamZ4tXl/aWnd0wAMImDQHFztBGo/h6rytd5fK5t5aDMk929yW
n9uTvNzkj31S/PBWUEoAPEIp4hde2ttDjqhT3D1SXMPSGxAOj8vtMG9OWfI5kXXty7Gh2YCBsts9
MhSurcEG2OsZ7Z3RKlQQnQAx+x/RaaBtw1pai6Ha2YaIELUSMkc1/TjJ/4QQWxqjj1LV81lpPWX9
dc0J7UiRbRHtX0XVDyO06+wnGCtL4EJVwhxxztPNgWJhsUa8Ij5pU+7TgGIB1Zd9JLHqc1oiDCJ9
pK7uNhqcrrWDg8qeizpfE36pdo4Z5mRDYq8Lm0GHELkRABqSbiLd7DxIJ69trwrJdU0vDTVgCJV0
lbZItAuLZAUOOugjOpPVIlxHFj9o4CjjbKUjVEKA9Jy2g3v0gGP8CER46AR5nHZt6emIgeZ6Q23a
y83JqIAjD0F14eETt1x3rXyUdAuMi1r23PvDLWKiGzSl9dlqbjHMw7LSmDhRrXjftN+DFhdETplO
ZVmTXQQSdFX2j2kHPFc5ySdASiyOsGtX9Q3jfSykJtMqQ7uKWWlChJk1REaTlYWVl2nC3t786ull
ZS18Ng2ciWH29eTiVCIs4N5OjiVoTDP/kua0ln8BNkpc+isDyelYoTI8tr+3YBp9cSXbn7GppRRm
lAu6KF3HB7qy3MZjdQzpQPpUDeAFIIFWNK0ifsGFReFI2T/ExvRAZ2xOr0Ox3kg1TzUg5jKP19ab
ZSX3xnXEqin5aofxtsCqqye2/bbwLzGIp9jzfXp/mHhQcBcFbnYJQG1dX8SuK5+pcrVN+Nb4zyxr
qPRGvk9REvDv6pf1n3sfChmPm+bBsKP5cW0ok1x4TpIbvBAShNuSm0v2FCnSpdYMKRY80lBqOEo3
DL0TGLh37gEiliO9IiAAG044WiCgwar0hvH1P3V/q07OdlCckbmsEt2LE2iDl64AoJCilgHCfUOT
/1gYT9miv4xEujdSF7iP11bqxaAHGbEzYLzprBYfZY7p8EcKAwH0fUYqIC/DA+NekLPljHd1F+5p
TgAK/YJKg0//JN1Qvce7J3+oMrla6JCR899Qjf9oVD7Z+/CMZiUjypuJi20cHYo6QCayFtml1/uf
bNqaCEG31nGLSB6RJ9+BYJlQIkgN2/WQGPz45ZTVGlXCCoYsPpDvDUVR8XEHOzT9Xg3HasgeZ8XM
bdsWvgG1I3QOFq0jyqWxld9ZMXEKtlib8T9egj4PslSMX5SajTlLtPG/445Di+nMxAQD+qwAJ4wU
1OQUa9IwOBW8kJxGYE4qR7J0BSnnVAb0puaJdvTPy55im5zGAp7g9hwpI3H0865j9Qgu5b3r0HlZ
LKa488W/ItjUjk1M9VNBvBBK0c6iR4lUIsoxHTDR7o6ftIvTnEUqktV255+OitpVGTNaSuJO6qkK
fVQUPqvEqhCDCNazmv4xRjZYV4MieiFCo/kZdJEw6lhS5U7Anv4CDfuBJi1nQFet1xx2qyNvCz3J
t0kOrUhQkwBF2VxsoZYrpK0Umxcb8aqbKeNFHlUdHNAICqSvJs5pzWCQTmErGHgUoA0lxZeKBk6l
c5H4/DKWqo0Y9LWwIl9qlA2IjtXhqyy85vD+wJpIYPo/sbbs8F3LXe/pP5l5NeokeYTi+qepCWUD
3Lath5vWl5m7wKhP6w+rdXjXHOaXOTAQemrOyRJews5MQVoazCLyqsioRbNcYrNcavKEy7wAKpr3
aUIZMAXaKHBU2WJqxPr/X0oT4K7Q53s1P7EZBvj+GEuO7PVPQ5SHqvIj7JBKIpkYf4ur7aJFA4YB
RhQgSdeaf2y+HGDP0WXDvxub8DTGj0KlrTe2WLWLxUxZLDPDMdnJ+TKcz1QnuOIUOIXUFKNTCh4/
e4OCPRK4m059TWKLIefgN4hEhcTtHzWyPpGtfsNSCagD/QdH3u8cv7/ax4B3UyqFZf72d9jn4zs2
d2bmhKj3QO5061OHjAlH5eKQmViFA/h3bum+k20OsScMhcVlKgGagN5P3ezznaxu/gjAoEy7mnlP
kqbiRgcCO4+SqBsXYG+JDrPeF7MwjNRumaz46ZSAMMivNvC/rquQNgAvI9Vqonbyy7NiosuEjs9j
cp1nfKTDTMfaZrnmhwh2KuH71Si5RLnOBxdrcjOfsRRs94+Eod7hVmTtHtchK0LUzGw10AdHWg/a
yUM8gi+j1WNbrGp6bTqEP6qWufv8EqRAivDPlINe5zy1wZQht8aLrpl5n2Au9S7iU1gAP9dU3lHT
A0m9PWL/ApJRjp6Vd13D7dKatFwBzdWU4UjVOR2GkXVxPQOa7pxCdF07nCeApj9yTwT00Car0bgO
qzO3rKxb3zVBmvxOc/JFN16HaJrriZxYFkJ2pmC3U5UbSoOcy11yFqfq8e64j17pZwhHI8nJVQIc
eZJzY67weVfRgokFy+ma/1yfM/wcji+ZVr52SnOyWPh5mDEjlMqUHlw2Zm1DLw6hFtrwJirapQa9
cdfgGYlCbIKT3ZXu5J9PE0YdINbB8OvKsLvtubayTBVwTIt7UFQaeF0Bwa06RqAsBPBM+olWDSmW
+qO6LAUu3tx2Aq/0d9gMFeRtpSfLx9HvmeNwWymTzsWsoAP++xTvBf2WCOWXPnPmFTExz8SehxJY
OHumjXj5TqWsZMSGxJDyz6H3QxBJaJT7nJW7mUvL7Ex3wEIbJptvC13KLH4jgPz6pmmgewaLs7hO
qki4ZZDlGz44EssFVgFZvRdB2Yty8YBqMWHRoDw9WDvt375RLJzjhxYMFO6fC7bjgpHSpxzdhAbE
H6iRfqMk5ozMo4wors8MZMasO4aK0w4KDzy4sDogQ2h9CP6j7S9VupqUx5UEM1YieOqEAV6xnKvo
Sdl060wtk+8VFiKi+drvQxnG+QVMwoUTfBeeqGSmZ/lHaL923An8D9/mxMAFQy1mSyfcBaoqZo0t
t0P+KqUNRBUcnl2Yf390kgUGz9Ibch+OmHylc6CoD9Je8x+R/k4UDe//tFs84qDEEGnR3mx1nQwp
6+s4KCx3aXK6yyxpFPqDRfWCfehxsKTjQH53/rw1AlgLwVPiVceF5ZDTGikE+GxVKr7vryqP8T8j
Ca8rDA6QWJy8hL3XaJ+CJnxDUdJdfOhfsXPFDXkGfx4XDnEQfbneUGWNuct3hNpkHfsQrC9RgrYn
9hSW7MEaMzO2eDYS7ATD/3Pn8mBzREocYEyCwxf5uEgNsTCEllNmSS2nVjMk5xPIQrqCfZZqah2g
jlncBCACqS1s3SzisfNy/9wBn0ysy9Vh0YFqInKS5380ZCoe+ULEzJYuwoZk75atDxK/VEm+O0j/
txFro2KKgey+jigXj6ygtlaXgcxycc0KulAIY3uJCd9YYmBvIxraOlpSe/rWqGF4j2T7EzIXrEEA
Qx5DBuZbmnwvqC8x/VoKRLLQ1w64aPw1ZXSw7dy+coP6JQyVPdKrsFvpCbIrYucY91soZoUqtpUz
bdotRzl95lg5i2Ob2p48EPPRkSQ9aNv9xy0JE1/vc9aKVTwAvCZ3WogkwP5ztRbJK+f0VlXfNZiG
5aFHwkxW2XIxZz4PSzUmdKp5faiDl1qZm5hzv2hnznmFkCVnr7Y1yg2vxB9Y8V0WO0G3jmQxLDUa
YspfvGFWMPdxn/cSveLtxiePCs+M+ZINHEQi5UkHOKEXnWEQG+pLQH9/sKbe3GXz/x5nGynQlFUG
2dfZriXWNXi/+hpTD9FW/c1Xv4pTBXNGU7+sfABqfpuNgX/bLabGtu1nv5BNdd7cZtdXlnRkHOyu
DJr60BM0XZOVKbeacoqRFa8JoOSvBrpnM3Q3joN2/nDqlBdUXk/1mM6kf2Gm3ypdaC6ZrILtDHux
lqlS+on3hVBSmsgYmk4NSYJNCMZIfOUw8IU/lTeM53wgObGpHkhQtF31wT8BWYo9i9818Aav4hye
DBYMb/TyCW0F3TIKB9HO5gLD3ujwsew3Mr8FYCGD3ryc9U+BLmj7YaVamrmjih/imnXdt27gxTmk
PhUQX09DLJ6LHRf8FkTaHL6rcBmGo/cbdADiW+jr2F9xA3UM0+b+VUlq0ILBYnQ6nhQHihiS+B97
+DczYYgs6CvxBv9NVXBw2GB/S/0OzWfpkayYhZd99ivDGqyVak9pHMHA7w7BigeWJgdJEMG+u/YN
kiPCUgCjsIDBEBDZ7cQ+AuqdJGqCKTe/vvqS3ylG6Lv8fcmwaTCJk5cmRIeoIAaQvP4dZG7wy+/B
xaQQZ9tWkU4C927ACm6EydjeZ9lh+u1UB/k0ncamAJ8RN/QsI4j3Bf/CVBy8UFVi/6zlANMC7984
5fbZ2DgS7qip6CjG6u50W/NKSmrmNNLsnSzCzMZGri5Y3nphjSPwMIwLeWso0najFuAgAy0ZTTor
OCjoaAWSMf6AOCMJa7RPLYvyJWfgCmUwOEMLt5JX02Z7UvC2AyA5QTlLDc+19NDoUuOzThPDierh
FUd++9Hk6CnKyybexwGkPwYowiPMGCC3e6MQ9Vmue9BpVR3FCgQlXGKq0tftAgDxZkljUEXmbvZ3
EHEeSYOUAw03lO8oqUE8BqL8RqfzEHrWONiYbCs47pkEtpnR4kExktZT+UaP/fd6RuVXiXLh4OGw
gZbnw9HOYen/hhQ1m4EomKXtZmkLWbY9OORAdrI2jbfLT5aN2iyG+n3BjqAq5nF8LSnxhxV0wA3H
AoGZRHfxzD5WTgzXA0a4ZoQYguJ00q5lSI3p08deHVDSSr6r4PHSEOxMifffuk8O3o9+/ortovcI
AltDzVY9tiGuF8jJ0vbt5E64WXgwokXbRcxK14nXOSFviojCZjFP+spe6gmx7Ht/DFdL2a2mRC+y
9ni9o9DgB1N5GVoMLXdcOaG5ZAs2+GWOhttAGtNhmVZPFs2uPi66dz+I/G4rhYURhteOZ65aXByy
aBBfGdNtK7+1sYgXcSSyiqwgHOMHdPTjsONBWMtO37jopp69qCzEOq7jkR5Y9nzHgFXb1PUmJOl9
nCB4jA4LDDFhVuv68x9lgarRRjEdnwkOKXqj8N5MC/Ghxlh1c5dyqVSgfueKuogYXgYR5FxT7Y6M
CWdgTGfL/4YyRxB6ufwucVKB5+5C1aYZxuJ1Iw/niTq7M8yxdVdBdfk6ndSf8vCNnQFvLk321Bir
KItDNp9AgCEhpnwlmCdwDxGgrF00xLGaSos6IF1TujR8ZrhSP4j8WueO6hk8RXoOIjz7kWEfS5a4
9mtK9O/lyss7LtD7DKFp5ToCj3vruxOnSpBL8p8REO7o53Y4AkQR35b6oIWUNgHQmzgS9bFNxjGF
pZfbyFSpEwGQZdvCXkOcDpKNcHiw5Ua7vnzz6qywuogiRGvqPP16EIKE1Ek8jIp1jA0N4a9hF6DY
Pa13J72Ucf0iWwcihXDuB5s1VrENqsEudNKBsnMH1s0Rnna7DAldMj1w+g5OAf61nJ7DN0PDDKYz
/vU/RK5tNsWxx7XKDcIy0c6IHVrhPcWKcfc6xeNEcfBGWvROUlsfrKHVkVNfq3OczFWFNGyQ4vYN
hHhFJlA5Cn+Sa3WSd24vpJdcT+GtfdPKiqXZT5bWxuE1VnaV+MOaNQFriJrBj3U2Pz8g0mlHzne5
6MqyHHLRR5Ca2wKQrYEF/AU98itUKNl6ue8Lxt1VPairyxqX6CwqHM9VEVHcUnVkiPBy1+w8GE4M
zCPgbB7etVLEsk4kBjWMEIvrINrO8UIG38urj6XjbpS1kV45rNGIn+y9mxBk2LpK20ecZs0W75p0
tAKtgrOYfK3TvqgWYN9Oy0NcR56E7faBRHlPmko0HEbKTFxoQ+Hp8A34r4tf6tqYyYFiHUPW2jB6
ReWfeyZB06XHumeKiIXXnsaQwOyrLSljlXtECNjWHrN2NchPsAnCAwy80ohrOofgGwgICIlN5h06
8JKNy2uLD7ynQce/5uG+x7jpjQ4qEHhGRNGgUHJcymR7ydkO85p4JnnMN5p6wuHgTv4fhAK6ORfF
hlAhIhxuWCRa21ilKo7Knj+YA5KLUtRZ7T8L4KJGRTMtVcV+lDCmqsYjIJowk2CFES5OAcw48WCI
kJYqj862Z+KUZ94/Qk/OX3be57OeV3cPsnYdvGepD59jx5mX9wt64iTc+jdIHdRRx+dAmw9JS3hb
VRGPtDOTV/1x1x22ZaTDxRJRezwqrqjN/fE6RxQmMiwqByvN0TXT8RKPMzbBsPcjjmg6hLNEm31f
/R1ywOhkfGDaGi9wkpTypFYXCPyUJdYMQZ4ddiyz6YpGO/ftj712GO9ic45j0OGt1qI9xbf68O9q
o+RrAl1KpW/+ztNPz3lTI7BQro1X16m/cSYFng0wUsqo/FBLfIoAnFBYHk9cnFBFP1G0Y69pFddl
MLqz8jU6D14RgQiAXI4qPGs0EwB63fSLqsrpV3prFkj5YSXD1JOKTdDP1PF7ZXo5fv9TUgJa3Rx+
CQb4owMn9f6A3P/gGQoRo8q4fD0bOPIRjNm3OWAqsNMCIxNU9Ge3ZTzCdmFrQ1rxpvCrXJj5uxaK
n5irGAUiGr2frfFjxiZPJSoEfmlYFzIXxkKiO1WoFJfUYBVpkjcIBPTo8cnICMJ8PL0CsIj3dMnO
6NSTbdI5m5pYrGitjyGKunqskonhfwXrelcmZ5mku0z04Z4cXA+ttPj0qw1I9SOqOFgpzO/lpeJj
W/Bb+6EcCxz2GKPWsjfEyAPi7AXecVuc1+QXioRr+zNZQ2l9nAve2qnNPuviC4m/0pjwNxrcrVUy
JLeWNeNs0v0heKijNyDh439wGEFFA6T/Ks1fZIgvfTZNubKeiAxMQjq9Ij/SAVcjH6qDgu7kHFH0
pnPddGlrCZ4JQTt9ULb6W+A005cHtKmhE/bSiiuAAHumujQksNAHIzKK4chxi7HW4Ow9J4lq4CoR
ZJIMRF6ax2zS7+ukNYoOwBjI20yfXRajzr8JTOWal4hXJby060SgrtjJq+L3jPSAdQLnwG7fDTRs
QNt+OWbxuaEmROa8Ue0RECFNOKz6IPzzKzGPgSJMdjWGW4jZZ0QeH1oTxLMdBSsJ//BsjkvXu0xc
p5w0DE7RAcioBn0iKD+3cJJhCLR7j61ffnJNKW/Va1d1sMwdomP/5BRuNw4ppnDPDY3cbwSPlAhI
3al9rggJ/8slLLyjVCYaA650vY+Pd/1EcpIfIlL1FXKESFSYUYMvXvYVxjegL+32PHCgydgIh2wx
DLCx6W99x1Cx6nYLbpCIVe0B7rPYttorrwq3UEd1umsWCpmbD9TUuDUYuXHTd8MYsJe+GyM1DK8i
Ac5GNCAXWtctn7v2u4pIJ5rvxGtkBI8/wtdHPZz051V3DAxHU+xIzejJmrFQ/jNqk68GeX5mCm/h
c/DUHspIW/GCo6456oVmbu7e2i9hEMXiUx0hKW973zG2aZb/WEBpHfdlld/dAl5UYN0C12nTiZiJ
6bD+SlLIWhNIyQV810lunYfSw3TKGwK1KMeYlTefHbEMGBTMfXxxmKcD7YLMjNRNEp9aelElkKtd
nPdo9+baI8/Mhh31lwAWdLRdqEKk8xjo+rZbpUHHbyWgPF/TCdUFPvaQs3A+QRBZnkvfviOI319d
ytYdUmPJS29d7UoIdM6o/XFhcoVbcbJQKbz/ESSMqyaiLYWB2PeXzpueNKRjhWMS8wpjYjNba4sM
0eQZQ2DKIZMM25+cZ6sAWAZwZj4g0jCDk/krzN/z3aHrWx2CGuduS4A78dFz2GhnBise+It9nDtv
LiL4J9Qn9n7MAtXgDmQgY1gI+yxr+4QhAFJFCEarivZ+fQORD/U26kYeBsbbwrJNPdlxd4DyOAUK
LSUmzYMwFKqGJwiLLBFHCEC1KcLeYDJLULMmWIlVRTZtyZqSEgIhCIIdsZ6qPRnSxV3MWbPmnfu6
nB+/efBW8aJQ/uBJOXXEOOI1mOKPeAQkOH0/ma5jeJKcJB2lROniwYoBFsQjDeB3uNMc1yJYK+u+
xUjKD90qeq77jNiTND/9xcaom5E9szKf02yxEt4Ilr5+ebFKOvqTDNXVig/vU+FpQHV5qF26Q498
WbAIqyN8foq12bi3oiC+15lXoN7c4vp1TE/d2jmeolpUowKPX2dM8WRBV3gCt66nCPgkYBAnzNTd
jdk4lYoXTAINLhf4+kOiLkxGFf9GDNFumEulxywpZawy1uJvG0hNZVcbnhYPtwzOwGLZjdy7ycui
vPWS3TZhc/oANfV3rJugzsWdRi+aYFyjwZXo+fK7g4udrVfh2jhwHDM4BCju2FO8wh13OV6/WgJ8
jPukdMZW78WOFwLspb69e5+7uwNYkLkH65turRUIoCD2Kh8SqM9XfO21+PAnPDYLcpqJzWhJPeZa
9fflzT60vaPmoCHeZR54wDJydwZ4cHxF/S7nyE2VEO17NAYzs+QbXnuziuwr4XqCm3KoSblha+cc
VF0CTJqQ1EpQ1cam8+EpowLqhJCfGPA8MTeEd0L0vWSEglkFMX3efLuE4Tv9DP8qcWgNsso5zu0R
NcsLW9ZX1jHae4AovjVhLfj2xXHPusK9IRQXvcJvr86XVcjN8h+MC7YOXCzYi+QYVkOxdtjZX2gT
lEYAefftRq5e/q83UCbTMLZH5hnuZ9VMWWoQ+dJ6WQsthL9YKWfaQhPdWtzZlx0IV8qJXHT+XNo1
VbbvLXj13X6gAXBNhuAi0GE9IdcLHq9YIWvUiV43XLk/5JI2zsV+fWfBOOpF5Sbgbg0blKDayVYt
s8BVm1iSXZJYJCwQI+ea0NVXm7v3r3auE3HpDI+xuDWG1sYg/ODNQ51ic2toBwJVQSqtIkRyxaZP
GrMM4rZlMZTpR2wUYGSzLZSHCzOZGuL22zhSuWlQnAcf6m7hIdlTbEKw+3T2Qvel4zhCo0/svNFi
O85Wr7/As0iMBUDAjvGkNHuUlgpC+TJH/8l57Tzqzx55P07/UObhGAP86R1y36cgoQxrCA7JH5Jc
BZquDAfu1F5BJ6m7Jy+ZY46g94zisrp8dpm6Di60x3Pad67XlacGObRLyuvJWFWBbJJfijQc6TRL
zQ0L2lajl/6nDKg4fK+/L44Y29yeYqcKtcyvb64DG18yHTqQAWqnwAusU/ddNo4A0WeJ182lVMzh
8YAPCDuAlXVvYRcz39R4Pkj2t1z/pkzeJq0OPy5EqMtMpi9SjkExoOdEd8Vyw9DKOpoVp7SQG3Ex
QYlVYsZLFL830Hc6DiVqgsVtXMiPRfrEQ796DW4nB/RC76cVs1sZHJrEa7EmSMDYycxOQFgGiEsi
+lfOu8T+kF3tfcS9uxReG98ICB18E/a7/ijM/T1S+Qe9+bjt6z9a0/TBIuNQCzLlaFT0OpGv6weE
u2k1bHA/2uQn9ReL8/nt1iyQtYZbc2JlqDhkXw7vsXQb5B5wMntpNtLXfiwC5y+YPdJilBVSz3v1
qhdxQLI9sFimERor1goRKsLrM0ZB/DRzCll/2LJEvRIWUEWNFplYOOKP64rRfbtSumHhQsGeP41M
qKqIgN40asQ07+kj93AL5jlfOl9ubPj/CVOwwhKZOWVE7m2Iu4HRPQD/D+DocNCusdHQa3DnymVB
AtY0he+xhe7pVKLUT5HE3WDzQBUinGmv2neBeAVmh1nUztLwI9CYtewxaJEt0xwNzGZKcjtrAwX+
XkWo2jnOKtFYjfLfN/JGoTCs1Fy8YPO4GdDr046/YLmLv5EJsSZwA/hOhICfSRmX76gCJhN0YFnC
Ehwu0DseK9Q6dpI0IIxw8HxpFwNltUhpPf/uy0cdkhZRELcDJ8Ojr8lcMX0B9EubfLy3ko4x4y9f
osJQNko4RqvzkChpB59yypOtxPotBkr+Petek6L2poDKE/CjpM+G1VjxQr/JyrFBHp6fblfenbc/
eTI9t4fN+qYs0kgBf3hJfj07rRPqLe7ltGe/Ofpnw48cr/3aIYCxVGps9i7cLh3WAonVctiopu68
VaxRwtwGJptpRP+bjL6CcsrBG/fahqG/stlDMWcl5NBQUkrhowgZLTXRbbfoAfKIaGbzB0Y34HxG
2JGEOZXH6NTc2FoeUu6YPFk7z9lwYMcnmr4oYSKkswpHwuiqE+CPuJPrILp7ov5SQF4iC97zha+s
PpiWUHS1qG6G/yWw5EmqcbqIlnL8HxdU5RWrIkBS+uVAt0epT5cq8jXFsG6zIHSpjaCL6pCT/41I
NVBbETjmpxLV/x0Mev2/sIooPLW4ObhUKI/i8enCfu/M5M6whp44qlMlhaz+0Nv3mOzuaby/f8kf
vhWv/BO0VoaetkR4SvksblEv5o8t1b3jsekjFniCUoEhlGY/PYaRVtncD4XmAWjNSa5leVN+sUl7
PJ40DxX9f3qKe46htOYSZ746Iz/gepSfANX7ntkKQE5TxfQ4L9acNTNgQl3pbmgkdG9hH5o+kJFa
NK0AKGb6WAX7459QqM8VYkdj89qF0Bar9BPis4ENY170MdKAiw3XeS/K9Pag7RtPlSHzqknQYJRt
ngKWgAxSgFW57+iOYZXJz3Sa1FG0EaJKuzzxQlqsmeVM7LctuqxxAybSobDgKqoMHSGyVJ+D0iQP
Iqk2bzVNYuvCAJ7QAU1sICZokprcBtCfOVllBxCNcJpuxHNEnjCwrgwzhyBcqizpvx9GtETuLe59
1mgipo8/xlypnfx/npAXJnF58RPe39u/zg3ESy/XbxzruaaMdKLjqifC+01MqS7eBV9xrHSt0nd6
t3f7iEE6LBBf6e9yjhrjSHpFEa8WFJW0YoBBjNh0yaCzS25E+Smn5zA5p2EFp5DV+w0/unoyDNou
AlSlvcMRfhgMvgiOpzbcs5Om3y+h/ZiTRTIBC1CI/TXqW06uOnBiHUq3dABag3L8poNm+V7V8Ssi
C4ulYjKeFEMDusHSYxaffmjRfhIlcfjozw+Emlr+4S/Sya1hA2XUwbP510lLnWy5NLY0ADiNmEAE
Y8RWCg8rHGXhPNarg1PhJrKSU6Rl+A8A4dnhBXKnKlcbqvKGd6XyHAkqpShCweqdcwiH+20Zqqo9
Ya3AHMNYMu9dPlEl41I6LKfFaDSDoQ2Wz5KHIB2LL7b3PLlgDPJAmi3ptKwwdJ1rFDYB2EoE/eXg
GZcF+/DAiFbxNuHalTJIms9TcfDc03sCO2NN+UJqr/FGFObPVuwmy8ZZuRbDBD4vKYQLp10wX+mU
4DuZ0sXZn64zruBYv4zcbbOY8EtdisnXSM+cE/UbWnNz7FGHZ+MJ5cU6028Ul59RC0E8aO07Pba3
MD7UIjm0BZCZ7b/huYGf8FW1wAXjY0WCwe9TLzPXbytGzkMIY8qawDshrP1Qan8Fq3KZSd6WpRj0
mELF1hE9WrRxlh8eWFT53vDLY6Yo4I9rp9weA3cWc+YD2SXyQOYSGrQ/+7+xLFnDo2AgUz7YAdYa
iFceS+vroXLVUABCh1bx2sReJWAFbxsNCIH1aaBA3zkRmxtu/xAd6BKW/PmEfmiCYK0zqQmgUzhw
mpJJxRH02FVAnCko4/ufHPC04tXJgw01bC32kjx3k/fUM0kvffi3w0yO21HMMGEp2QtaKgf/I00L
bhp0lBkEX3LQJnjOoOkaYIiVXkzPvRRs3YxURxT28tuGjDv944TK2GmX+atvjZU0/Jt0ygeJEcHv
KBH2KF183grYZ8lOtU0c8snaLeowC0/Gr2sLhWjGCdlinsXL+zinp9UWzRQGLrrcbEGI5DKiBMKL
tDRxUeinXDrZ+FlJ5BLV7axoZzzRCu3r9eEfacxlXDpjqwA7sZI7p6ga20x+y3do7nwES7o9Bnt7
yEuUrfmwtPTlWbRZ20cOaNog7eP+rAeYy65MnjWhCwtmyxJk+5fqjVAFpVcco4HTlDiSoqrmew/f
DmJ0pI1iicjLJgxzGpGP6U2IVnwPreNsddkNpOLPYptw1jiWyYDNX+FhqirpN4nbT7TDr+8Wbha3
oAfMx0lnOTQIJ6PshLJCYYZP/rP4HjcdBWg2S44c4CTi4fKIwxJU146kHp5/jGqLZLYDsB7Kk7F5
F3e3caW0Vys2RV7hFZShRogdm5lKhzFU5KePpzVwkheN7dJk8ajGTwvOpyjdOnq3T7GjTsdfyOdZ
aApEDhBtEr8JlSxNjapdmneIoCBCFcA8H+dBzlXEZ/hZJTdPSvQWWpN1hTy5dV3Vi8WxddJigpbx
xhe8laMHPFqnSvj0vSokPRWVvvf2iIuX1lKgz8WnNZlbsDe+xrEVkYC+BT7t6EodxCRKHLJR2T/y
lnA4rNWVinrTOO98bjHpRhSbetXCQ+JgF2wzRhZacoP72amTXurWJnzGYMA0PuxDD79MiCwzCaIH
vMi5aR0uBwQ3nruvJKWGkS3c4FI16szTXFLQuHHHmButqacLkFCt+0o17ClCDKCXGHMJpMkpR9Lt
cQ1F6LAvSXEmD94shZSS2dotMi4aa8cZNJeNjUBw1c+KOVsn+cNqgVwgkfDp+An2gBqlhvPg961W
FiWliRZ1640PzpM7FfC2f8yX+OBOdRzHAuY7KDe5xJ+nl9TEQK7lDqo512bLttc7NguLtenGX1AW
E+1v/CE807h/uON0/5v6+2X0u8A1Ws3e9S0zfUc2GxBcpNkSDbCQu1q5qfByhb/aSimnrsM4bSqt
ibYHVPYmmKdeOOx3YrtdqZlosoZ+hX3sUzTbmmSp1fUmwqoYVBPV+wpv9ACbPMmz8uEJpcx1wUyK
8cleiQCrdiT2mZPy1gEcF/pP6QK/Jn7ulUEaYrkSjTTio70I0PWv28tarvgJaPf3cz2PBz+AgsbT
mUyC+Vxce6I7uRqGK0v9FFg/tZvyrDFhJbZO3N/IS4/pGoqN76mFJKHMkROYAkcR0QT/7dsmIFUo
fnsforuTciMNqMlrPlXq1oq66jBNrnEgRToCB873D8jV3VMIt+lrZPqj6c06neJHLcmKe7SOQfG0
yRyqKC3XkkM5n9AfkyVcN7nEAk+9NujmJZj1m1cYsyjlJp+Yihz73b2K2ErIV2Fq76m1d4JhAIrX
C/Iq39B+gNxXIZFZQNb22i/eIa8hSTeRGBfBFcXVIlxiZmoWnU1fQzaj2+vNlQKIoXOA9rTK6PyU
oTiGxy5Pmg2qslZ3sykh8p46U0qmWXUMz7lsT5n8I3TzHYbZBgTaNaNqx7K4/geeMSCt+7PIGt3k
xBy2eN2FavJOcTgCxBpRdUaTme8tTXGMjVI0likPsqArmHceM8rWc5mBI8TYtuXVx7+mqtGQCz/M
VhoPoGs1a93RsZJd+adH0fyWWBLOTLalSTlu/jEz9xt343wymOD1jBJLsNVtxIxlQ0IsbxhHCmvL
SwtPomzA8TeTFkbc67BGBP5szAoCSlOQ0J/jrcTcS8vbquW2Gn8G/G+ZQxVbsg8T2wqBZk0R0ZWD
TOe9oosLrFH5a3VCSyhKQP6szg1l8sS85mhWXtuKPfAQa3EUhIUb3aXMuEL1xI4c1eXNG3MYOp8W
QuTER/14iO+piRVETwUFa69YiIZmJp43psH6pvmBNJS1AbDWP6GZ7cw/tS+DXofmt6TG05mnG6D/
6ey4hWTkpUrLxiBJgBHvHLCHz7oQXODpPvx+rICbZgv49/oSKCVFYw82oGf8AHGEHM1gBzbNSBoW
sGBwSBsEqREB74XP4wiNsVWjQYoe78nK6eJdG6D0puTKmpAfmqtFrr2NLdsavPI7AmKCcarFjGpN
Jdw9YDg8aBMQu7lkPh2bXu9I5zlXdY3OniMH+sRBxmKmiSrs6t6M2ac/rHbeRiAkwDxsnBTkWY7l
aS2KyJOKVsO+qQhyehSP243ieQfkXNMZLuHJx4DgXKAM97OuOT9GBYdmFcCV1Jt3linXtTxGzPca
5exyFOxQHBzSjbCvqbXnRreBYKlLxiIVgG3uysW7aSzAj0wk2wN70GMCxNDhsmK8slMbOzR3jUB8
5y5Oeq6ApBPyuPENZ4pdDVUii0VT2gp+LLp9PNbYzJx7pLF80pqfibIwjUM+miN8y1b2toGBrnvj
G6KH5zFN2xEcSUx3TeCw8rSXcQN7abA+5vxB3jkSissEnPOG/Fq/QR9WtoB+oEtTsqS/Qdf1mjxc
UUwlYES0/SlD4/Z/aAfoKyWxskm8P/x97Kq6odaXFEM4G2GHF1WJkdhHC/vYo7G9SFrbTL1Y3J2j
0ANovp1PxAPQNDrZSjSBhwYbeOk+H9hx3KQ77eGeXYuryVRnyCar1pDXgXXM1+JC0bg6UOsuD0WU
PPgSkx2ozr6ScUSMIrrPZZcgmyykXNSG46U80fPHQNJNe8sZLAQx+1eMPe8eYUgfmcRZE6W/gcXm
+yVJBul7YXhGyIDeAvYvHo3pQl9MA4ydV5AT2d5HDuh7Azd6tP9KoW7M69D+kPeHT3nu3ux1RmoL
KOZZA3/eAyz36XkR7LpIs6l8k77exWHbN1L0AVWnyvZOnf2uKTS0Pjmq8I7iC+oXOjYnI8XA7GJd
rCL+KZuJ3yf93303tsVjlCmgaakqWMw43URrzTdTnIBpd1U/4sd1P9NoFKn8UcleJBqTxfqg8pXx
71tfxIMlBRn9pI89P8DWlAZZU9SlJFzTI7um4VJrlhcgZXaJfuPWDP3Hd83I979EQ/kI+x69A0Zx
CjTsevq58lDYijvJt3KDdxOq9DEHYHau7H41uvHygo1m434UfW+il4hcvJD+jkaDWnQ9Ngqvdnnj
qpaPBCBIkidZvMf5CuXObeCysKVAu2LCGjjL93LBh1USmr+1A3AUYiD4mGGrmlRIdNKP2JnwVLxJ
DHblajQjThpCP2gxShzydbiEpJRJSID7N7ZVtkBlEK6D1IVMqKJ0gm2ug1NdCHkmOm7zbdmAMmCz
7Lybgy9Y8dHBw9jD/uKsVhejmVsQXovAQQx5H2bIwjQOncXNsaUzaqBQJWJCNGn68AWgTFQRSrWi
TQQavjZtuAZ5iJNYvbTfCJEWM2/6zbo02SXgd9Mo77yegbxNdcOHmvPCZhMT4BZDhH1jysfrqdtF
kiXlKLI5bm5/mOcnVHUQhZQ6GcwuJRB1RJ0XTfH4S5bUkyGr6WGdDggwkLtTkKwbzYcbpxSQorrr
+962hDYHMeZKzg0vIhPEl48V4tOBt3wofn+p0URESHRzFYtgmd7bbZQ+Xsac6ZE+0i0QuLYipYWW
h4z+pQrQGVb09wvSk5q3Q7va3n3IOdG9RJg+k4/lVLqdHpHDyBC2jtWXgVAPDJ2liaN4qQ8HCCTc
lz8pUBlX/rdhWNwYHiWM64ZNlB+1S5UwJV74HEAS1M+4Ln/Eu30CA4l7BHdFz6gaG1yqFp5VipEu
NLoPhCoLtLTbqu9iio4aF6r+VB0UUJrtqu+UjtOdVLiOueg+LDAqqCTNb0Ln9hjOLRfU87eTrake
3MVbyuv4yVcLuIBF2l4RVpNWokCyDiFP7TwDO7yfIQ2itrbPhSAx1PTlizI6UfbpjmsukmZQCuO+
/ldWg/n/O3uSOsaU5mQ4tYabTpWhA8OqeJ7Lqa92ejyjqujN6PoPtP2B2aubYGlYEhgT4V9QhTFg
C8Ta7n/QiVo/A9LvOF0AKdvt7sew7UOIVcW/gdVKjvvHHjmIFMeaUhXNDx02ykke4T5NgQo+hGCF
/jyr7vKT0Pr8rWh3+qKkLF5fu/J0hhbGLjSuEwC9v9fzb+Y6RV8iJVIVXaHQ2RtBMxw7tNpmXZxd
b+szT5eyqJY0T86uzUu4KqYn0F7CdqYNA4kxuA7gJ0peSANolOVe5AAVaeaPlbFJbUrD1QaqlgIv
TMTqozGmnaPBWfMyceLocZtg/hX7zm3NquYg8VdqmIhVm1GKLPJfBXR6JzzQWBhCSsuonwu+3gjX
WZau/rkaza0+Bd+oAr02JpYmLc0KpWZtdtXmAHx4t746rFE1WUu9zKRKO+Dr5k5tOjUlPKCDyVNl
ZMlZ7SrPqhBGh1HtsmZJyZPTPr35sTnGJMcvuIcjGTyRfE0Hl63fL9BTndc4vjh9WLMyPYByx3on
xPbh5cLtIGv6v0mEWTYjtCVIraQOxC2u1D/OGCL2RXqvlQ0OUmM353VWf3KNaHYjM27Rmo7JSIoK
dSRCPINNhwz55H5JSJMWuydQlGQ42roVnHvqo+8j7PkR7kE24scKEqwrEDzoxmfh6tI2Lo72U62M
nA7zvfT5QJmF+O+EJeCAzQtft4djCHPRSRyeO7A9KduMKZtHq7qSSv/vHu0TTKxuXYvDX7Zi3O+y
ur6Cp7EaGu2VrE3N/T6mTW15E/qjsTXg8SD9nAHD/QgRYZ4ywI+YlQ/3ypZvaR5QiLBB1+k7ZV+R
hxrz6BPC1zB424ieju9YNPsAZ/4rTqCSns9bjvor46Za4E/OdSw/ZlEO1zOSNaxTKnIX8o7wYmEU
+lq6lYoqoxtN2Jd2yUniS7Q76tg9Thf+5/EdtCWh4sFYotN+Pf0DM1ixOy9iK/XJfDI66DqN9lBR
AK7ZoZd0rVUMw5vVBr0B6YGG/vsgSsgyDemZgq58LankRxzlVfAvUdS57vimy61Hg7aPSEuHWBCN
b5TymUKq0a2RyehkiU9nAI9qpEtOIN6vfgJuYA3BtJQbxo58f9ZjQHPJU8zhuQReuA2rx5y6o/4h
tmw2cDXqp28pMxcDDCAgn8FQW5RhRsDZgtOuD+s0CftpB0a9/8MfcqM/rfl+pqKRxnMXBWVR8jqm
1OQlHyPsYipNVl9LHu5nFOXczc99olkNa69xUw0Imirj6ReHW7hCc9OIwYMiZkvWM++7GaBllVYm
N1jBqfdRSuRAzfknrLhQvTQZRF2t75x4kxLVL7VJzChtOgikvN/B/wQXsWmjUmtIQQIf1ZineLev
wCH2Ku0NJlUFiAGCbo+YNITACXf2hHRGIpYcIEpdJwQZKTo/o3+7idh7W7rMpcGZD0JLrUvijHBO
bV0bKuIRQmSGGRr71Rk/PqoA42uvJZKGuGmcvdEkxHPuGT3mD5SCS3TGMIvSLPNV6hM5fKsfUxnQ
7yKtRKIhSELXMhRCDSiEbTYLLRUTv2pj5kmrXrIzTJv+ZNEFo/D+1I8bNp2IwSQEFZW4Mn7+TjyS
OclEgrEW6Ii6GOiGlMnSUxMZgePKHPhvTXF3NlEIWU/9lRozYkH8nNIerFGUJwq81/AqNtk+xKi0
KoDEo7BkIqS0+D15kdpq3ink4ytbM3zMZDCaq7X1mChR0um/uhFHnmwGFQSGQKhxQZnBzQmcDNBR
LqLjN8CpSRXqsdlSI2q3zFNjg7GfXNkMjvc0ok6ZPVMACsDBHtqNNhK+j03Z8ZEXrAzJPtsOtzCN
+glhzXqFdv8i+4DhWtvwVaUJWf4MabdXwI4fLyNQI8HnAKFe6Izusxf8/0ADi9Wce62VZmJxh0s9
j/Jtk12+8apbEqAR2qygJhiQyAaW7X86J/9Y4R2xyXDvi1H53F9hOeLS+e+LfpsiWzg0IShY+HeI
/l0jyTXOautUq8SclUZALtrR6TGuGF8Moy718/jyLg0ovZsThFxPTWBhnSHR+871BZ5r/d6oypoi
/qWVbUGezh4oQAL0wTWeGiSZPeWTpHtFv5FQ30erI79mbbT/vYwXMeVYm5tFIPczQ7TCR79wuexM
CFkA62VRv4HQ/j9tE7DwPFeOfVMPsu75+JkRL9cYOvDUiiTG8gRTRnIvlBjFL9pamHZWIc9Cu/Tt
cCGxyd8RLOIEr0u/II9qYb4+nDYop4KGU8ELtIF1zcV+od829pZD88xRSWlFduuT9oPft34bvZam
D7f1hKY+1mqAyY90BomeBLkk7QvqFyL6ovBxl5O5iEJuNhELnKd9LWJWwmu/ygo5RrNqE0qTKEhM
vzkCIZqY7kw3u/Kx62FXRJyNbs0f3yAAufCVF7wkJze7amjDNu70cTZFaneVI9kUmb5+ICCOXHP+
/ip3qGAdHBXkmNtWFva7mzukxuLURNGFOTP5zWzQXOoavNl2ByZ29g98jbvdfsLT5FME+KIocgvt
nillGtz0MRFyeedY3/MIz9yJagyEOOQv/ai8njYXF/QLLU5nSAoI9c/FEbPBKXsfNNntvDjNk5fV
JVpnSkqT4UPPtuqq7GuH6S1E/GmNVDX9A63zl9M6q6Rx3hW6NjT+W2FuGMSFDWsShoYKinYyzqKY
dm8RwL3oykYHzOusjh0vxB814HBOgQP8NofEcwvT1DMHtjknkovdoM1QFKPxvFYnnpoYr/wo4OSI
Aw4rvln873lKW1kw4uuyyvY+Q+QrdmYbo/ia/ec8ivmk6YLye29EamP5vZnr2gMWu445Gxr2UacS
CDFp7tnsykLg3WHYM3OvayxLagxpCar1x7Rk8gGAin4745MVT6jGqpUiDhbdHZZsyS85GhAiUyMh
+U9/TQsqaCpuKiJVagbYYfm6KPVKXZJChx3Dwr2751ZQg8jkbUa5zqy0qeC+4CsYKhns35dj8t1D
HQSGD6z6pMtGHiY/r6FDKKzsRml34zptAPkREagK+K+vF+wJTb8qMky3p9RGKoHbYg2+L8C4D7nh
XVQD6kMb4fsp5aDwV1Jx0Au8dOqyz3fiJ7WKQPwZzFj9YNBvPe4HUZZqOkmZZW2Y8WYI3KoG4j8m
m7DodR5m/iCMZFaVF7uOqH6msPQhiMSdxfga8MlVC4vJ+54X2x289YCXYwACDh6uUURdpCL4ltSn
vTOo56HWgpsunleraLk7d3+uIRb+4BwWr0BpR/gDVn5qG57Miz36uYQGOqU5a5tv4yPdm4JZqWLz
mK96sXNtTgPto7RhFpSLGDfU/Pj1Tr5qgXlftNtLc+BvixzeWf5czhNGItSlILGFAoq1drJoN4NH
LuhGKo5VO1hx9m11+8PjZuL1po+z0ELMgQmEFzSq3qKne1hd1Wtx5who3BUjQBYziXl8cyaXU/ps
hkkG4sEO3YSQff5Kndd+cuDTtexyfLeibOlhX8ByI10UkfdauE2qo47Y6ieHATdO5tIn8x0MK+JS
Bsm+H1piK5ja93Nsr3AEHOvH04Lxi1cg2cFlKzEonQiLil7RhiyvAibPKUozR1A/X+MCy6MJaWOw
N/OV+dceBOMB7nkSW0XSjU0OG4+A2KGXsHMjHTSk8BBUze5TxIkUg5/NJMEVEpn9hgGSNuGTWbGT
biUNRp8o51ttcLC/rg3YjLKZ5RlWWrqFGF6oUZ8t48PEtOKy36waeDGyfHDsUoOktZyORKAuoNqi
YYZlNA3Is3U2EJ6zrfZbkF0+tOVbxM6NdT3/F5BIqyoXC3d4eYsAxIniASzVV5213R3J/BbS2fRi
tonewKR2AXM4q9ow99YnZ/i0qDbPyEbw0Mcf8Z8ouQieDOaDwyL9Zs0iLasCkLipKyZBUXgbyz5V
XWujo9ZNvTqgQ3cg65IyBc4HA6V6ZYDBAWvkf/FnP/CqSb/gXx9b3w3/fMxJi8wlUeRnCWt1urC/
w0GFKcCLnHEF9WWPfySgTYQWm7kwS9GbuI2gIE+0qAIFynAFzbzyw2nhf/gbyxWJMjCrjf+Cg2+K
mk2K9OIava0OxuOdvgdXeXbZD9h+F3nASwqGjmi22OKCIC1qjZxWEbQgHn6eCmakYQ/mmURLjBdy
s/H3zqIyxexsSFTXc3+FIENCQQ21Cy5AypT0O5fqFieuGEuizqd9Lz2ZRYKn4kKBg08kPXvUIgIs
q4rmn2K1sHQSj0GWRfhZu9gwjbef31Yu0oR/xNDG6rpyvlWRNo1hIs1Ui9UOcWNtVKsALBbOds0r
PzQi9MDT5NH4nkFrunabI/0xWbil0TYQhuGOj52mMJ4ettCukYKWPdtIgjp1jBXLjYdodfgi5ZWQ
KqcOSyipf5Rxm1/K77zhB0HmPHUUwUn6SGJ3xNg7W/bN9HmDCqw/qr4462zrZ6HQqX/f/LFL8lqd
KlSpH7JRjRQy9/TSzj1CKwdf7dRozFcMljFfopdfIpSrBytXmb3iHJfpVUe9QtYAu1dsjJr3wokU
fcPAG5mRYt7MBPkVqtFFkRueJNUAqkEohKZDFCA2DMrNNMuUqen8uILXGpkxnPj9u9JE/uaYih33
+OBfqSr+AlhY9mEnG9ruGpsM7S/0ZHQjI2GBdh2rST1NQZBrz8ceHWiPeJJhOtKLZquSjiff92zW
Kqo9GtTM1SknJOzxg/rMVUsEHExOcUcSkOgCK/lJgsDnKGb/V9iFTtL0dV90c3LtvxlHcAvA0beX
y892+81ugy9xNT7FABhmNJBj/oOtbrzRiAsv3emnevvhBeufqzzTxa6HPS0mi8aNBnB5qyvhS10g
aOC4q5HgTpcPCRFoBfzguKN1vg86JP/zIeTFobOKn+6GjWLDKg2PJQ38dLm2ls+d+1nTEG6rJXa+
ijjM+FVR8I+iEtDLVvBRFD04CMMTGbqHy8dxt7isIasTmujOlSWu/CFGdyJJQu0x7eIHDcVrKHoI
BYnmh3Fk1w8Bd8OOn4Wy5oiqaQY/45xNo/idKeIjsqMZlbt57B/QXPcNQjqJBweLPES573ymnG74
zgkAnqI7vH1u3DwB3eNGqhCiC37A+A9BQgD/AIiPMKMoOXMae/pu5H07V3lIcjwGRSd/BwBYVSeF
pPaOJ+6Bgo4Q3L/qgVynzk9yRbpJqmvwWOj8HGWzH+x5xsXZUfEV/dCLDW3zGQ93FGwsdYrcIXe9
BWVuOdRVeRBqanQcZHvExKQeSMA9b1HViNELgUWG/xYLL0oSeofxr1PPGG37P6UXOivNVTuXBzqa
o0BQ32JkB2lRpEssThWDjqHJCNrPtG/ozbNw7s4EY1iQIB7037/QQ6Px7ZSHY9KyBZzGDYiWVj3F
V2CGsUdQHsfA9OYZ+H+J66LYaGy0BChEwz8SwXLZ/Vbaq1tNBGSJLLYAYMBPAinNQvn8UImQ/3oz
atogH/4s4AFfRQPtEL16Avj1SUsQRLsQwCFMhY0XOnVVH2o2OTv6KFkLssKr5I+f0WlScH73hVC3
BqTARcT6pQYKjx6NU8q6ZEVYjKtY6TAMOxvF14YFLdFE8HfsvgR8jZaxKCyowkLj71j7QXkVC/ap
VkM7C8+7qZuR1GUXn3ROiU85FsOVA3GtuzaZ8V2lUGOnZC6tUBTp4oaCZ1PZkv4uv7Mpcu0xBa4z
dMh1EiUg0EcDKlSuZKhQ7xcbD4iUB9d1Hjqs+UxXnKjVPLqNWkQc1VRQ52eeQ+5fYqmZ1kbeIJ/o
FHVkLf4nW8IyF9T8vIA3oYPW90/zpx52WPIK48Ff9ix5fnIiL/ruUbZMUj8Sm76HSwBjjVDGqKZ2
X9F7SFyehIOWcI6xlWYZtpq1BouPIWmKNmfpGByEU2PQcm321BwV4yCLk5fcAuoLB37wpKLj9i6o
a9XkQjkbBI/zSKxkCom5/9p9zIP91Gps7061gcmBY7xMnXRco1s7fnXqffHZHIiIB3/KkVe3Ixd6
VmRy70Zl+82sEOgYudMI5zajmc+hUGZD6q70+HxyOebrCz90Ogn9AtlRTYDpsNt7rBieuBI8v4W1
Uzj5PUVfZKVHF02uMcEtSSpMOJnkRbUru2eMbo2D3GvndKc2fJKB+mbCCgYy53PtZ30Dsjt/GWwR
tosddQySrTa5JlNU4kXeEru1kisWyJ6HAAdOaJ1rrYGRpVRJkj4kzXkxL4WqkAlIQBim1n1Bwfwl
qU073vdr1GCriRzQC8S92j92yLRWHViI0C1skWy4BxHxq9WAZWbs7y/AL2qOKK8qvM4DE8EP2yCs
R4NN9anHXazTro4vcrq+ln5ksw1zBhq1kOZcjrOqBK8ZakA3ahQwh0REX08IVJs2ir3KHb6sr4QO
9q7BnHi/3D6w0zNMFglRQYGtDPRVfePjv1hwYIMcSJ/+FBc+PtMqmBhHjyW3N3/aN6rsqabm8R9v
BDi487iTNfUrc0k39SxIVxorzw+c0r0G12v7g5VWm/EcIehlXTUICnC8tH4CnGxaTIccOFRDTmc5
uKc8/a9nYBpxZBKLtejyE96rEnwfixvvqVTdmqgyQmIuvWkH3Xgm5HjpAm2ZWh8LMvvL6gGVQDcb
41CZKE+ZRvVixtRH1XmjWt98mab7N0IkHB90/uDylAFK04tWZjFa8dJAI39w9Qzff3wI/SWVOxgl
5ZMxW3VsxsQXU7oL6XXd0PRnFAd/ZD7w95MSrkvz+cSES02CLc7uIjAUHC5dMFFPwgOB0MeBgj3s
1cl7x/uRCPVKImAJJ0CjGtDwGub6EDShGG+LwyUS0JRUSAZOblwkF4+yD/PSJ9BNryTVJFDngYy4
P1iHUwStTtnWiuKSHcwHSWfhEC6C+0HIC5FOij2jerDDKhtzY4Ky6NPPz2tkwJ2JJ5zBDge9f4Cg
3nTCJNpDOMCENZlFUChMQwMU+sEBbnxM0QeDcBiDUE/XevBacMS+DWwLhV4QCpWHsgixaZpn0oFW
deQgiPV6Gdj6EqUI3nDeaCk6zy9doO1nYMXLG881Il0hs2QPJuqbQ7YXm/B/mptS3knB/1m17DPQ
E0rDJBE3U5pXRAtPV+RWV9w9zH4qQ2xFtCPTlSmg7WGei8UTp0UVc8FE4aqSMB8g7TQhmZXE1oZD
e62etORCGrfnxcwkLYEAlJukGf6JJN5M3uEglZTgi8X6/KaPpQKJx3wIldXJxOyhjO/Efw893xxW
0bf7uLpAcQVPtr+PtUN0FYwYMtrRGl+YW4XB5cJfdLq8h+e7fKJLbR/s7FAI865t4R+bEkyOiHzS
FaJ2YLXA1+Rxq2dEcsuO/u8CFX/oGMmXfNVegg0HrzX8EfieGqo4iisqM/zEk8+srgB7esC6LJo9
Op/DK4XPe/P3x1f2KGtx7+pQlo7/VZItIzVWbvsKhxWIWIi7JlAiYahef6APDPoy8i53PqafQsyP
zFWGqHof0/5mIRGh2MjbWAzR9MhJmIokHLJKp2kyn2jO4EMoiIp1AI6dFLebKg0+qczx3mjw5/yt
rx0XqyMcIFKaZz9SifcuOOlfrdAh7G/8zbjsBocvUylda0oosTHyNCje25vSjMBfNQq3x6xx7bpM
3ZMgbFUvTi894oTXqM9Abzw/63LeAo1pKCYeJ2DGVXdocGPJ8559cUhDPE3Owb5119YFYSdklldE
jzT+W0mcsfNjdRPRF7xrbvnX4HAVSD+LCsCnnIoIdvtxDqWWKu2LCfmG7AuiuEtnkN5qj9nhZXEa
iqqRMDg2HHG3TjSkuWoakgH9Cq4bZwEf4ZtLQF3wRMYOQns7mVSysGEi/jYHBPfPluZnMtiIxKsQ
bCfvEQnaOzwwL++3QIt8HoB2JPr+SZte0SAkV9RUyi3Lgv+FWkWTM/BqvkqF2pWcQJiM42UidlKn
uLfR9Fo9k59wKuQwXee3H8z9J6wgOyDydi6KZ8HFjQT5NSEylPw1tt20g+eDq3cNEkpgRRaZ8EsE
dXRExlDTzCZ0ZnW3hgD+vK2dzR/7jES/uKkx1zM7iZtJxEPCfpK35nn2r011FZV+2DxL11z1mRKw
RAin8rWEUtvFV2aUgO7FCHTBQMWhiJVsFJW7IDZibOSJLcLJkK69N7vVYpH0oCKdJIwJ9KIxcxdr
RSMxEBirbtZ1oQZ49jNtN9p2mV7JdbboICCky8w7fgsN2Xv6/nN7Vw6axqVXbrSkQqKwg1s9o+db
CBfn62Y665pz7P6n1ihtFLb6eDCcmCbPlge3FI7ohmp1fnnJv41jms8YRk182Zg7lC1+yrXkhlPN
XzRIhiTGAmvcSM4mIyaw+vTCd67qmWbSgmSOGCIp6IsdZVWgoakMvmR88H2Fa0X0/Q/+x2g3bNHk
qoQCvL8WwGr/y2FLO/wdfGnvvhZwsCt7F4eIkfgL57qQGh7goc9IDylSBDnbukOSxfCdqUR+mNfE
2Wz6djRVUyPLKH6miFImybW1h/cgOwFgiX83d8jCXusV2yCyqVdt1M3m9Jv49nxvzU8xso2kez6z
idXkBg5b/jZc8cVgwfu31/nHv2jaNQqXdICTGTBxGLWkGYIaz1GMRoVa9VviaBnmKDHOp/ESJkYm
hJf2d5zWjYANQ0XfvWDrzgjWkDe6QGxZ1hP2jR1K9rfSlqf6/CRr72oeR5/L5V20BVRKHHIihu95
NI/p9CKqt6pKbI2oE64r6DpabYt/AbjxfyuCCtELAVE/aaQzgyFnPeXKBGGy7a8HKlRYWv3K+AHG
WgkDmosuPNp+5jJVhYMul+2rJXP3+xXFbzVOMEGWy71WuSiPm7T9vgjfyOCWrGAMmNTWMCJ47dJL
gTma8oc/uVZ7VufzL3qmvS2zfBVf6LoUciHllgLQMeDaktAo0ocRhE+rDV+/Mb9REJILr6BS0oFl
vQ2LLpZIsQTp/yjDCoNsuZTcN7V4RL14f7Su8apGl53O87d0QTCzk22GjBPjhM2+KwjZc5eG9kNu
7asIDrgPiUy31XC3ER3/duv12JmByNp/NXO7ellNDwCN41aGUh9btTYFkrfmA2GTwm8njiqGfwrt
VspMreUbEdDp/VahQzoMzOjQ9UqK+kr2EiIk99uwfhzKXK2wfptQ0IrESy/ELCCgQ1phkjnDygPM
H4Nf2NvjXMAvf2HscNVd6Tki9ahD0f/FR8M+R75h6ssTHBfxzqX1ZoKD2EzIxDHgDVXvN94gRSpy
zC2CbldWaek2Ql1OrN6roOk4BSktasT/MFNUKI0HnbN6rRsWLmiAnUAUsTPjdw3G8QyxPfh6owiU
nWFGSl3Y3aJxqS/VWb8bc9eHkfmakiGl5a3TWPH0CuU7E1ShUOGRlIRgjZzV+XDeVh6KhcW9moST
+slIngzc4Tyxk4r6oy84CulhFrYgzJYr7OdMKnb9lJNQ1BSidlB85/AhAtpPnzM1bYTJa432I8WT
tUfUzyunKBaOcTuIShsRIpClNPVN+YbQOj+eLR+nXWlEA1LvxjBPTl904eocjblw3r4ztgxTWeDd
5EM+JxaNFpSfggDv+W7eXIs3Dk7/qvH6EJo1Jxq5p/OIrBBSoCQQME1Rb3WQH0e981SPxZIaClrS
1rqB/eomLDG8xyWV529gSPAcZUV+ckSV9QzFkbAQW2JaZBvIhA6o1BSurEzZDot5Qde03meg3b3z
vOOUCz9pMzyiZmD9gRiJNPUXab7mM0SREVGgWEjaFjj46Cr7tca+QKc/b8bq6tlhp9+dQvvVSZMf
po/ykBzcUHzl0cgMAe6cym1xBTIiySCeOtcI9w98brcdlZsS9EYpG21gd/iODj7svSOgzWJuM5no
ngfvnFIqfPPPP9xdg/K4+L8jGuUGYD8g9vrCzqTDvwBypRrTh5VoFw0kpj+17orHC8XUZC6GIWjN
vjIQReW3FJYFCsPzGYk9+C665DaI5Sd88NSJV73OBuMwQUb5GgHULRTIGkl+yJoIM5+VuaI1bbxf
YGunz6mvFGpT9KVMeMpDCqsLlxHWTUxf8c7hkNxPmWxhpXtqwBtUtF4pK5/N9Yma5n2Xy9YSZ+y+
vH/rAFKq4xZOrf4Ck8uJS62fceidW+i0E5cbQ//rw8fcB4Nl1me5PKJjiwPC7w6GxSaWknkfpMiz
ukoWaVhsB45WtUHx7ca7uFOy+1wP0iknHqPJQXmI06CdjQ+8x9tpev/8Pm16IIbuSAp1VKLYyerq
9sb/Sp3YG47IYtmfdBxQ4FBHLbS91amaxGsj408F8IjMmk7eXKUXQvia2JGK+vSDBLgT41+BZzhY
ZD8vu7yomp11eW5beZeeHamEuFYVLfQqq7zdD3r51fzryJ+CZ1m0weaoY8H6CwiVOISIHmb+cgPT
ogsTtyqOnjH7QZgyR1bdETtOf25hQafEnApKYDVEntWS/OH2RYLBq1tlXp2yKvuwnHCDv+Zvi6OJ
pv+aH9LL8aULdWpDuwlMZs2ykigE46iC5VjAm4ebqAc219G4CmROwVi46+K3zSDGW+TgpoorwcEw
z0cQXxkTnBXLGnzE93GaPsxeH5ZCizqt6HlmV8SCvaXAOwGVt97HJmhJHc5zqE0Pku9DzkVhKQbl
SsFa2Weg+FOjdjx44FgqdWajWen1nv9kV/J4W+MYyACHRl9Ha8GVPGBlRs0So131BaB2xuJjzyil
QbK5M6qZm33ypFyiVZGSB9vRVHXDVB+NKL/gfW9L5n4Sm/VkkrI563PQqyKwgOyXZerBLQoi5FtE
APEhOEas4iH34g6+QtbGTFLgTYba0DOnjYmvIqN5SB6xjNMXwVByJm1VcFDglUw2wNnzzFsKckpl
0NsqHgMDLcVYgp03Z5aG78v/VC+L2GXtjMpkGtZW/3w5R4/R5jXvD7FSi31QBzFMmnFXz5RSUtQ+
W00yIntc26LjfY+cE96MXL2oCb/t9R+sC3fM14zp4b/bO6ffL3j59HEuGIJaVD99V5oLm/fYYoPp
O6sET151cxdiUOZ8804S+dZWQk0g9T0HOi/hj4rU9VGsfgExuMjTEc+AIPJ7ej9xceWR4MBiN7LM
d4RuxeRRVf41ZKUPD/MJvV1zYZRjFkY/kZq11bf/01Eg7SUWPTnhDhPT1rd2+XtV/xcxdfKKqty6
/91asIRi8En884ZdNyH93AVOSeK5HKpEAGcIExzhG1xDUzEsMPy4+4q32I7hXBin9TX9nQCx0vIv
2hqxvLO0qH8CedRJIFki+wg6Vg0Pm3/gk6cDEScHXEW66SYnm4jLBK3pTosaa5tXCTqi6EpSJiVv
R2C9YWmNveu62XKFTQ/HEndtNrRAopgJ+cGUm/RCFK85pnXPISbwjYSUG/pi+/mICBYiTDiyQxI5
83kz2hu3+0wOddYCgWBtQJKdYNK7ySKtYaF2DVPEeRFvlLChgpf+37vIMPRJCSftLVT5TwFs1+YR
67Zzaxpqoa1vj57AEsJhcGV0nvdefLejDdr38yLrHggCdAw6osXQAJzZdraf1TH7okyB66m4hdXD
R7YlU16rGfDxtkkK3GCpEvGPJXNLsAL5XXV3pGpO4QAZOhMlfh0V9je1S1ZfPddDvlkRdYLw4FaD
MqX+Hi41aIV2bEJ22G5cX3+JyDr7lFaO76zS32Ek4+4/ikftXRf20wdPeLVNxBplZEtf7h6bzIDo
kCmQMfZN/yhlVctkDvX9q9boJ47SpUEAIgE9W5Th5FulQCmZxkRzJ8Q/lYpVADpvLj8l7vid2fDg
FpqOrhZ1ewO2YnKVrn+InlJ0+/mtKzz5Sc3HuR26/aE0Cr+qiRKnCSSRuG3XdE7FlIh2xIx8lJ8A
xyiPEFNjZudod5Hh4WWNwecoILdCYT9ZkqbUOqJiF5TmlK822yBG/VE+4EwkjbFWoXa70N6rzfUX
go0R2UcyWwo2soyAB+sKDrpW3ETr7BONvK+G26gaaHiWLDw5KvXZkdpAq8EvHNJuDWELPeytoL4y
pk1U6cPSc6+QDrLuq8d06bLZokhbQ5dzwgb74GcI18ihZ8qcGr9/zRxTgtQRZQbQ9VzfcGPRN1p9
ZcqRrthTWQToumTVmLrqpnoXs2Cbux3whfAUOK03+meJvTlGf/FicJtxZUnn+LGLIKffzs6OKNVi
QlA9fYgsDjLm1f60SXXPjFMUpMJ6dpg/qOgCCloUn5iLIXYPqqAAPbrONNz52c8YLLRumaniwN4t
pIz6o/0DyRoa98xRRkDT5WkK0Q8GqSOw571STdnARqST6dFsviaFP1dDoUcDgay4Piyvh6N15AxS
2jmp+ZWbDHtWmaLa5omjdbM4Bqv9nk1L2hz8x2qH3xWo8dKPW4ZwYck5+lsC+dh+ufLQJcwUWOKu
4O2RkFI7OTM3kMS3vOzgsT4ZQismIaUwrprpxXLYOXwF2rxNy8kJCtBV5tpR07G7T5872lsb36xG
SAcZn2RZamtb8sRjS/Z6JSdanDmqLvw8ZPx8JKnahK8bvhtarTbw5bQB7vZWgsOQoDVKI/Pehlnu
6Vr8z3XmOFYvCX4YgbaeVx9t+OrNqMnSxvJf5VTTpCgjIDbfysgEO4QiKOPdEz5loMcOxiVaCVAZ
6XrFAuXLpmmiNVUxrwpAAJHpYdkeEnid24h0+E45Hryg8wxyqwGE68V5uhExztVKWZ8QBrh7kMgQ
FyvFLKJ15CmvU2uEsQ3WFyVgDiqfwTGRopNU6CgX2gqdn1kBN44wkNBzc+7kg/FGMvp3/wRcFUDg
+hLmo0ORG/l6ykklBqFxOlLjq3qODk7Lgj15pmiSV5sppGSxwC/ddrQdzOnE8S0PsK9CBXmfisI2
yJWyUP/phAmS7BCeFxQY59pmk+ydKIT2Pk7XPKTulWIvho2yDiXRjhYxOcjYZoaCUECmKNo32ANO
d38LlIJDNacMhJHHCIUP0hnukRb1TYn+5E7k3CWoGAHoQxeDYVGiEuR7LoblpKMb4MezgGpODt7+
SVVXREQrNg1TAf7Cr2w2IcgqmLVrhm6CEvxwKEtfQTBCFcOD6qiGpai4pOVMcoEBsPn5PwbWfqIa
UZo20lhTYS9D34qtEoVi5viXT1lf4of9pWhZizqv8XkQaLmWgOtMmjVRy3/iu26Brn9Zuzszyadp
zoizrNJKauc6NXKWj+QTMsT3G1nOwFI6yvf4JFuADH5Vu5ewh0zmSQtR6CIrnGWQRqWe64D40yZl
ufKjq0RmL/41fmjQ+lplvZ6HddY5nVMRTlpvDEliZmMSNYBX18BwQoeqasg6ATWagwAXglNN9XS9
txXUL+QkI9xmZED2kGofALnwxKVLJxC+z7D0UYKVH0lwBDoDKQ5dNxg1SKIpIT7eF8H1bmmji6D5
SC9Q1dDhD3wCM4j21MxzypnIn7DBooy6JG0qe9VxZ4sE30r3eB2YcBJf5nfnZdjHYSKDLmCac7Om
5Z9n333PJchS/AjSikTtbVk6LQaun7c6payCvapv/865oHagOjjz4M5ffkECY6EjaFLifEoFXb9J
eYbvgOqchrIG7nzMwZahOZ0D0utCO9dzo8hbpO7ACtFdVmKgX7GByA5a/tIzE99x61eiCifpG2ek
WFBMi2430vFqAcKUf04kCNNbnoWyl6PPPFfUEVYly+M9iLIjgyqSj2aJK9SpJezofCnYH3oFI7hE
WcD97C/e8vkzGjcHHrmXBfIB/T+4y3vztSGzgPlodmXfXoKD3s5hDRLGDGjdHoJG8i00L8Yb938o
uBmjNXKkcBxHNWkoOIOUDdkTSb2BMYcFjXvfdgpFyXmJ00SpWjjrKewHVJZdJSn4adjeIYLd5t04
XgGLmRiCUwrW0VFnyRz5Z4M6B7e4wy+SUQliU9H1Mn5svTL1tQ6KgBCeb9OpafKoYhgzkyv+fjcv
gTGGD7dWQIruUi2Pxi9v4KEfxFKEo10BuH9Lpv3JOcQqOKtN3P1afPhIqqBKxUsVnizVx4HwMY2b
9ME1THB9qUw5fGPd71RXrVmUvqESogG2X4MO1ThhsiI6eSEMZmlIRij7d2pcCDQVjwyl2XVAOIzx
g+2t92HLgd2tOrbXLs8w5NEKQTSK0TC1pbtiecfC7+1/VE5keBEkairftd93xivACzK9We0i3Qdd
qtfilSc9diDihdkZQ46o7VLmX5mEyQgmQIZBZ2wdBN2LeXxeW6TcGMDftwBjna8S/ngzPVHpl0lG
RaaAIgWJ0O+ydH4B8NI+aTcNdgSfXN8FZ+4+l5dCtmgyzv+22DdUzvJ7bruIctNwrrlGArJEnmvZ
KMsCqvM85H2sEI/ttUKnJMG9SBWpFrC0QQ1m8QlrlOXQzB1v+/aSyHwgrkzDWtQ53Gjw1JUuKaAe
zUZbf2cHz4ijsDDN+HfRO8NWAIdi6tVi7FYYcarhwQ1uKKvExqwwL6IpMpTupTSZX+yH10n97dN2
gmnz+jLOpdcNhPlf51IL1xRRHJxqjehXEVVYOO2OsBvOZ9L4jMZBKYlNsoXJx/3j7b3lgThUTTms
9r0sRVmV7vPGI4J3Ix0jYlqKmmeu+kT/VGBtgQMVUT5FGN7FRB/8clUroNAx2wUIBfHR8ldF7GqJ
I+i/2NyNGHc/3Yw6GU+1g0dMx09r1g+S2/VbOgsTZhzjcsi4YJZH7WotdX3cohQeUwhacDXwQUHE
CkXPOzJY3eHtXoDRcsytlzDB47xZTHhrN1oeyfMlyboxICJEk5Z8dmpn0v9Mfh/VjbmGgVHNmZYI
FNDc9m4RddsLa+5P3+7sVwvFoahPYPWx0uBHkkV3xcuA2z8ksqHn0vTqq3iU3Pu7a6Vw3A48sNUb
FWvG9mvaRipBZT3+x4fpQv8C0ud/EFQYDs9lQ12QamuA0vsqSHfnde/Uo3E4PHaXE2x/jKXYNxLl
jZcGaFP7No2fL4BlNtOF2iuceCOIuyo6t3Sf73HCg/ekjZnABl+P0WZ28cSqOqWzUEx49TGErErR
nw8Z7+YqgBTT50dthchf9IUKyjW8q3n8qPCMd+ngdcSxaURyIkwka3r7HuQvkALRHNj1Hm8Yt1mb
BZWRWRA9P/ovFsDhISMhYmFoDomKyfZn1//IkUahB0MCDBHHJyRWkGN/LvWHQC57rArgrLug6LZS
nbi1t7WOziwMaZAXxnsguWP+ikZAiyD39He9VgooAP1PdLITOvn9BZXdpqdtx3syfX+2Fy8ldPTT
H9Rs7g7oNANKdh/qtkSIFPYob22LWMdANEADvzB058ZzdnINHixVE+tIZksqrnPQEQqaT1EpZK23
lz2arC97fkOlHYH0kUvtviwYQqyVbsdVAzyXbgAKQSS2gxIChzkyx0nO5zdqt/xLAq9wIGeD2n8F
sqsqa5MNn5RQBItYbXxxpfnmJSJqTKE9dAfjjBEy015mMSdm+tAlxfBCFLSAek5XK/vUEStlGONj
LF0nizVAJofD1E1TSDWyD45/L1OGUD64VQFlEW19Y/iDv9SngVwaLvzWpAR0GR0fhXD3fHPAo2rv
UvO7Zvbv2nW5VfPS6qqZxQuUXYMcgj+AHqb8Qmc0x0G/aSNf7tEaD49Z7xxint8Z/FBUrTeeKQLw
HXlboZbu2Yl09ihxBRK6Z4FfPKTavzTaB3W9psDBuXCOcHM2DpLon0ZUyNwGapyGsO87DPvVZnVj
rZ1njNY29xNtfGwZtrG5pE4oWge72nVOriIIlt+VRjegHtsZ8iVXZkQ88NCGDMe6RTsUhucnTF1z
9tgeRpOpHBrdAz8wMgnndhdVUjWXl3g2adQy7welxOGdpBmr4Ny7h7Vyxyrp6HcyjbriQ0GivG3W
ncr0qx4rgVleJD4d+JbpQw5qbfDdIjCaNWu1fR2qHWhgOOYqMTfQhb5GnfYOxdPIBWWZ1CHQ6plj
KBVpyHoy6hrl/nEl4gKRjbZEzUbhkSq5ktOd2cOGmQVZLgoZs2e4rbf9/M9OouOBf7u59lV1sxho
0yCEbSdGEMV99+A/YByYIRxlo2kkHtiRru7jK0aYQdaKPWIOWJRxid5P78ja8rNJ8yXgzReO+Upr
UvH/Beua+/MCsFadAucr8Kg2sXBIwKTcRPshqFru7aUuWTLRG59I+w5wfmpHmwIVGZiBb+ObmsTt
VLqBIUeRxQAzs6S3gGhv376k59glIevo/SKEq5rst6PAiKMhUrmBA2ppiYfQY78pMZ9WErszt4/d
SqJLemuZ+Pa9mxQck+Lfg2d4tBitmvyhhbvF/TX7HM+hFZhxtVAF+AdRgmkgWNX63Va3ezcU4694
sm49PXb2jKdoL9vYCvfeB5LE1DR5Z6dJrVnpSDe8Qm1fSVNwyAnkoxJGIpyA5TkXoMtnIwsLegeK
kHhDHsqfyA/41dSxLsJ2RwL9RPgzPS2eMxGnrmqgSVxrVigL4Vy57mgLqdhMVgdzDMGDnMIDqujZ
wB0whnv25YOv/RaJzh1oAi/CqsdQuxRkj96owk+yptqJ7Oghmhq9tXqsHFTsbrQM/z4ZpigLbvCl
BQhbZgDb8yXmOVtkdWt6Q12CBVtIRUBCWg1oo0rEmGW/oAPcOi3vodTcya57xg276MM+0WYNdgLf
Jbyleb3GqJFwOrGeLMoA02gMK6ByKBKD/QRfhsskapLDDhwzLhyyjeVYm2IUQad40st+oUefztwI
kQF6EWqXGqV5Abz3hpJqcMDjLZF+4ICG0711hGrn9mtQGQS+fErwYhN/H+ybN27DrTZBBg4uvYXN
CLuaMDlJRg0ERGn977D7kWgItiTXNB9qVi58gVBcOmBLeVjJgMW89j9TCfcHVs8ztaU58eznFu3H
bTmsLuqae4IlF3bAt2LBQTVrT82yH+QLUxV/TBSABZNShzUbI3j6SUS2ychTf6AlUOr8wyAANfQi
084F6xv0gOhCC/rTXlSEcDZ3OkXrB3hLfgmW1vybhlkidrrgFzHylf7nun3RzXJme3EYazt/Jx2I
1j6si75alLoNqivwrTSTjPqSVQIHxabOsLvM0mka4A3o7yFCKAZqkiZHt87Mr6Q2Tb51FvDRtRbf
81xQd730VkKmqJgjtJj6LWvT4D1/XKXtuGt0MWiMcsWFLPiPJ2xdGx4bKTx+jSJbNMEKn6Wb7H/b
pWrIDc7wC6HrmFGPe+VnOXFCuDngD7rtcmjZ540oz4oTXts1ocaGZOgd8cTQb4bFYIN5Tto+zTzP
nz1IIknx/H+hvBoepVTnyjwyQJGS8ipe1S10BLPIslXUAwxf4bgPBrlt+ftaAWILv0NVpEKwu2NX
XugzFGSKb/zRNC9mDKHwWPaO+AxgBor7kIbO6NBi8n0oZGZ0cTZI4t/WKxxqwrZUHWtW3ssMpZwF
3O3M8zq/mYO8I1OnaWvj05Snma+fKgUJRRHoUqP3P9vzctPJez/qvYQbiHMgngsbWI0/wcrse/eQ
Ph7dIAXfREFCQ/dEAAn4aI+CMqiWFgQqOyrBLVqbahm3+X1ZQwyLmG7mJD4kr00kWnUQa7gK2YYX
1dwNOw/nTsZVKBw/VyYU02E1coPD/86V7P4fyrlSpyQOg64zVsXlP5oyHbmTa75gI8wjZQBny9YG
G9xD9aFd5T3mkXnW+L3nJqGuaNsc4UJfZrub7wM3tkd9QJ8Ek/T58bzbJJbrAhGxbcuNpuq3HNgB
kBzq7sVZizucWobl0SrFvHC97KVAdvkw//UzoSviDuplzTbxSEsob60IRC9GiRNsVeufospRfTio
OL0/gxjbdbJf93Svk0v7sI+U6sWYOJF9o6zL8VQRMwzNYGC0V56ULLQFfKYVjgpfS9Gov3DSbPSE
STHwAn7X2mMaiI1kmXmvygjj/Q0ftdd53t+bQoKhoPxBMpe7z4/Prg467GheaxO6NCDo/Nt/706V
B3uhPv7xLCBdhLh4JfOO7iTOlcm2PipEAJzaA39h1XhQX0MeN7+ByPIF2nZsgDOnUfU6jOjxr/zi
1MmvtDU5oV39Kfu1QWRHiCgMDwN89FNI2I0tR/kEEJ8RarxXFMlvllarrulZEnREzEqAfPFLL7j6
j8thMRVhnJGgS1s0YWRP74ti/FVpPtvowmQGE/V73rX9Lvye/mXE+jvRwyuKm5kyRbrZDT7Vgwl7
H4NblBX22vT7VB9wkccqV8VqD7uQ8FFvglgT9rFuW9meN10htYH9ieB6c0+PFEMRZ50Smz1PiqWJ
IvKOsyTeNiR4Meeo6PWWQFDd1/TQYvooSXT0diTPHEys0HCBdqDNRXiS2D35AAEHndiEpJPfv0JT
KBlFgbzu3Kq3kcd2fs5IC4akZRWWlhaEKqKaP7e9vE0IJBcylHbzOpAHll4+nOqFvGZDjkjgSNMG
0YU8SuHsgcQGQFYxpyVW0zA+eQmUXpur7FR7hLRBeuV9lxjKo6iZuigoDhw7TxXDreBQOmmo0sRL
+scDNTfxd3AUQlssC0j0MSpPHGBwFX8ouaDRprF+uASxV2R7yHjPxn3aiinhHs/raUQr8dgKukEA
1ZSYwyGdsoDQI6L0eIIqZ2SSCedoJ5bhB5dDNepENmxmUsKfP4AdWqUPR3IMGFE8De/1GOGIx7XZ
yHQo5N1+uhwil5GfRTtg9ppBEaPBccm0e6Fnzq7S8/xtEvYcuDSGUt9jsX+yIL/EGPvj0G3cpiOY
34jIN2VpRwhhJHpqlNGM2mqe/961rG8H76pVspZL2HjLYfUgRMbt6YWtO5URNUinlnOwWA98YuAI
SQe5HVCkX+nUrVb9kP1Se3un3IS2jGj113q631n3zoK3dytJ0PcvNt+VnbtjC2ZUoNmuGlSh6vRn
VrthfAO46+S3vjXd9/+HgtpHZRTuIgqshO91KPfvxNcdO7/dBEbA/lVBaOvbGwME9F5N7ef6AVw8
XxT9OcnQIHsrOCIKDTJ+tCJLmFPsBLzQ07sJ5eYOM/v6XftUFXQ4FdcaV/cu/+qKetdpENt5/7ju
8AlGF6LbXQQ4LEgdLb/YUKcz1xjXQKYLjZmsrOaPHCTVVakD/znSm4psXZgYuyGHoxrmAQ99xMPY
fF0sEZkGfDKdblRAw3xeitso9bsQQpGFLoF2jvOoF3PPZMqTL1v2TDI1xdJlruw/gLMFATdXu4x8
bVe5ETzbkTV25qTY1TtsTdA+WPZwQDSNwMcHHwR9OhjqcuEBwhLE54jt3c/4r5SLey9ZSoqJeKl4
d/lSzV16SIlv8npKYkAbPE3I9qHfZ8caG3yVZAi7UwFUiGfq4joAh9REQA3b/XjT9/bA4jLhtwVt
B/pgkUUMFbpoNCN9wYGF5fRbBu4+2JdYhkEEdSqSL8WN1940859J6wYMGFNeCu0PYzqxy7HjvFVV
q2SROUR0y0GRFr+QmHhGS5fV7Tt8bFLr93BwjL/dNuwmZ/j4DIoWwgdoXNYKlwKg3MBLvn85Rz1A
54QjAgM2jc3ZY5ulNAqaOkEz8ulBFxIt0jPXtbw6MMWxvJVxKfMcjDdl6MIuhJEhzmn4stSpxKLe
G8Pej6sKCdHleyIxuCfscajtRyuB2wGRylDlwrnGejoamP3bN+LKHXyPq3zg7COlS4KMcLrDn2IZ
PGWCgPqhraJbWyEzJ0Bq6hUFtT1HCzrnVU1nEy7fhd/WLxOoQOEmeCkR/iYg7Y5aOjNrJebDBdmS
XsWMR60OWyTzW2bWrDrcoQe0Yf3cFrTVSGnzU3PHUN2uJuo6rDhu9iuvhnF1AQot3TaKiK0e87aU
bODHIl49/ZqmKIZntgfjG69CfesQaW4zDrRZwpBZS8U2v9rPw5Izgr1o18tciCnK4tTXySAQqrKy
stHbvQjGwp6cGwVw2WBXpHOitoEElfLcAwNN7yHwzxGjnF2PQziBH3wUD9nhc+uO29MQUz6jAR/U
+10DbS0B3t2/4cxvbL8OxvLYO4Y0M8lC8dhErs+pArIsgcz78oS5dmPV3HNBbKTK7RHtZXLxJwZG
xgHjUBTirJv1FTqu4Xk65KN0TnHlldjirfQLoniyowVjpPfC7teNq5/WmZuwilYOFX2gwzw6rskw
25BbYsBODfMbs+B7Z2dZJB4z/38trSL10a4FwaPfZucT7YtVGazO7XJfD2ySxwBppUEndvuVqYh7
V1Ooz5ZNDWOMMG+yFZ/+a0+75/zPjmIAuvzu50ollQ9kzEwqpx8bLHt2fTuMdJMoJIJYPFaz6olw
oEvqsnjlIq/RfQ8JWCks5SC288IWsVKSCf1RGcErw71NrgmZIykTR3sxbq73GgyLB7RWHB4rc7Kz
yG+Te8dxSXQuiBPI0ivlgGZuItGOk30aWOS+sDrxnpSc9crDaFlX8oSmI7APRcoAXmD37VLdNTgG
Ms8fwMiqtWCQsnGxFoKWLhpKLvh+YKE8eJAzCtY53kMgHkjUGfyseSOo8VQ1JquFpAV7u0U1B31B
4Twm5VbBewzOvcxnlbZTgdjLttyPZUyO3VGi3xUgtonqRiYThm1La+mdsLxgVLkqXvBJf7hoKGqO
UVEiMk/qWc+3E/p/b5SdBp74P6GnyJjHFELJGxMd+VV4bN5W4VWS6etZE3tHWceyRIO7xueg3LeW
Oho0NVRwDQprKI3w4KFsf4DFcllVZ8U7/f4nhiGyRpsAnd83D+uZ2ApOSxF6sCUXBavmSwmeWzDe
n8qM1rUntOCMxz6O+G+IlnbwuCpuwUVF5+Jj3I0MfLLWz4U1NKgI6fr9P1/9ljZuOlBoGFG6wYNR
Xc3z5ZWBrkJ3+Np1biTXc4PvRRodimdwfRNWQBMkX8Sp+sv+z8UfNSEV8Cnuh1tIuvIj/p+MMgPz
YzFOWXvyoI9clmeTGeo8gPLxmdOk+9hUJFW4NDlDqtF63fwAxwBWtTvYMKA3LxEUU/OnfnuRMS8s
08Z0jKUEgpi5Oh2Gt0NhB0AQ9pUNNe8hMEXqIbin1xdpWDcApGLE43t/NytLfoAyP3AKuWHieHrq
eQusRtD4RvgJVUVIKQyBTMuGsJRkwIJsuCsl/DFufGSiapGU68yjNWdM602e7/dOBoWUCQ9TgbFa
edmfX2IIIAMgKZPxA13adleVhu0LkZ2e3/HYhnJQXk7SRR9M9fGF5hvrSZNpL2mv/1gTgJBQ911m
AeVHG0J20T4HfyI20V16G1WYBoLi43QxO9fRl+BsrKfCPelrLikRBzG7lkAXG10IvTkGBE55lL09
/txHgh2w87upQOVEAcfEl2aT9guXGUao1twsm1K5NlBBAQ/HBb5jkdXRtEW7z/Zjbevv3I3QFc+2
NQVJQpvUjj9xasDPLwQO1128hr3XYqpv9Gh64wkjGMTW2U+dpj18O9ZwLfA6Ne/zkgeX9jbGIila
YzIfHAjXE0EBw9GMeiLDG5SkELHJTUTHHFW4qduOpN4CFRjxYoL5hkna0UU9eqDOfnjCKIDP/yyP
CwJRhG9F/+sVNDa0JcU/TDNB9UgRPRHc+wUbcWMld8K2VEgfF8kIZQmLmHJz0Tt+gFlAMmIjCSa6
nMJn8zsVZK9fSSExjNL7/BbhaxCWVstUMnsz7NcvQTeO8z/wNc+SaNiQT9V6AHzpRjz/pGEqHq37
s0rphykpmKX87vYE/J4oa565fPNXJcTLEqdkUrhtBVkLc8SZfi3o99LHQWsWstylRVAXviWATpW9
rC3ejd8JWlAVb7cRZXM+i1TiHY0xkzbU0QuKdyV/JWb9UmfngX564i5sFhQ5g0JCrA5bFmhDD8jD
YwKzUpzMJTUclU7cNbSwllW/GEO6hOVW5H1etNbgu42g05ka4CnVPONNeWDTddlkpDoUZXoU1TGE
cDPRHObukdRK7lgBTgYj83Sd/3MwMqjzZzA4kaFZ55+SObIt1wvjzb1Y86LL9a6j1n5DvniaZRlR
15ta6blukNb8HhaV7mwUG56iMN70wBS/x4DivF/DOSF0OILh6UJ7XMvv/lVbmwJQS7CnJgME041B
x2jz8f0BjzQBWZLuyZFreN170I0p8J+m+8dg3ySKew24/z6imLZXcH5kGbTL+0K9sMdvg50nOUPi
Yt1swNszUSP4jaUi5mTFrbml90EPltY/fFbzuFkm6TZAoDHDrtx7/519qUYnAhzW51WvoBaBnytQ
NBWK7e78B6WRSUa4niorvoQVsgwtQY4+2FQ/f5qQHRSbS0xuMmZkIqipxE0/jXkYfPmizwctVS9w
2iz/4EQZx2NNFkaRGa/FtbMsMI1CwVuFAsZAAybB7SB1BH3FXnLM+AvKJJ/MVIkxuODSyjT7zNio
jWlu1F9FTIRl9hVdUDNBOuGLYRVZstNzyAFCHnJha8NUJReKazQmNf4TvV0Gg9BX4R8mlHmmtSjV
jSwyF50I5mrX3/wPYg4/CNzzZb8LK4Fyzi/au67JtyKw0/liI2WDtfFcm2d7ITEXLTb8WqYaWHs1
vfGUF2MBuJdOOPxuQGkdMLSSngvryPNETYdDuoQWZiTR9X7F9NdHZu2twhAn8i/805fC2hSKjZaP
aGFSQpWFbSkep4U0UFOx313itZw2A6frX9NSVAg0aJnv1tB1fKW9+LV9F5vWfbZENmvNdpspLPzQ
j9afO6YNXlkP8Xj1xsQ5jlBixd4l2sSdNJYuptM/8Cl8LlYCHjVyPky0rXmWeeP627xs3Uet2ddi
/ktlmHINFN6lO2tshkKzQCpk2bLICHoGPJb0l1XH+iaTHsOO03ECn7q6LvxaQYPUzvc/6pcN3vWP
50pIbZFSXboOhmV/Q+0Qi3JqNWIyV8Y7n7idjWGFluSrqFHbu++nGRX5px9x2NWtjbirCyPFmQjJ
EPOd7I5RdhmDp1HIia2Wc5Roq+c7CUs4pJJzMFFOntBC4kDige8SE1z/b7xDNG4KNZ9NeaR0WqJF
wIvS4Pw42WQzdvSLtRAulMqbq5RJHBllPdAxF1qGBsBX4SuPuNIla9O8NAsm+oJSPwpA6LKQH0uB
NPR4lbiL4BlXBv0BVuf8mZAADjpxDPWT8Ob7x5XLFc2iVFklsnqSjCAycbMRRFBTnWDOsgpBGXKu
aG3UXBm9XmzoaN8dDfSwEBogGbrHPkxkK93ESe2o8ch52SOGh2ARRZY/8H245IclO5SUD9x/arp9
zfSl6sWzzOw7Jp+EL2YDRGaxJKwBr3L7ayS8jmi8SNyb0dpvPn3CgOp+MMupI4MqswqiZWo+U0DD
9Ip3aaLW83jf0nkDAExggevbZw3t0V6Rt1ZJqXsetAj6r35cRagCgx+oClIatiQT2uMR43YrkIwm
n4ALewVnDJD9zlOTlnerQ35tp7nZ3G2Wp/vuquyWDalJwIJUa2YsBIQKvivBIrjXDu76FhGSsTeV
BywVT45owqkqfKjej8KHR5rcmJkT/HFaizwfhMeIeJPp6rXvnsf/6x2p04cnKN3yPG5iVnVcWISq
gkrv+CvK/RDju5dg7nC4q1arXJhC9PXA+iET0xgJyz8r0SdC5FBqPhZjUpy0GLHKb5kFNgZFladW
uYqCrSddCoN0AGmkN0YKtkA/RiC/R+SfXEFu0MTamPJMNBfoE4pIiQDCVOZR+y+/lkUrBQiXv/cs
Lv/fZiu2rHsFASBFbrgU56C1bDwcLrKmFU7mQye4QQu9UGayy+GjsdrmL2lRlFtjgdpXS+p/5nRK
UhafvUOooHT4B6GnCFrMXJekoDHW5SHNo9hyDaktN41wqbE91ZcGCsZZGUT74CZEXI8zZ+M/zu3o
sVazOtQ8Vk0q1dPBHDvFHSst9+AXxcyQWUi25YQ9mn/nyIi1MAjxekufqeESNT04RwmCXvmXZ/ie
sDKPUO/7dl3S5rwb7fLbUm+wmeHaypLWG90ysIuFYEUfkrhl64u4QkPR2oD9jUrQAiA1occ52MOg
ZIEWKhQsDw1ckykR5M0v+O+C6DJC1e6ulkZPZwfu19HXzgohEyzvM2s4SdSKlcnUK6ladmHZCgg2
E2nY1882+XMq/T3I4rAn22GuktoG793W4NrVvLK2KByDXUZWltz4guWw0Q5XykniTvx5vPCy1n5h
0NEG0jUjjizg/L08LFOH/dG2kXW1q93Tx4dh4+Snh7SGSHqfsJlwUgFtQmglt12nziruqqW2dF3H
ty+2bLu3Xz9Nm7adgk9baF6EUTcwyY6z4z1DIXUjOUhM01PiT9Cq9jeE2YEomaZdqHZnJC09W2PF
jDElRXGSt37bl8t5gPNz4khtd/RDUFcDEkIXyh4xmnCkFJejAiGzjFnwIu0iSvatdlTDT89ddBMB
zaZ7BR5N32pM3bNT4SDjpfucTTkXD0bT50+PO3fEX6xhXsuljn7zqtjactg8i9TJt3rsrim3Im0z
DdkBppBNQcFWKM06uc9hlSJae/4NOADU2txTof0WM1V9h11RSLBu9+49GRm/MkdcpOrSe0571zG7
x2VkxUpOrUtDTbsUi/7b3NQmgqu/5hg9w5blGy5g7S8zaiWxikytnrGsbX9sTZE4LZ/+dyg/8L6z
81FHk2GZgGOCBQ02mZ5NpcUefqxxlsQ0Gw4xu3VbayZR3hhIqo0hW53wbrDepX6y4AgusCpNCJ6/
OlxUpmlf6xDrNstIajYC33+C5f/5vM0CQTY8E01lurW6no/D88HU1Rc2VubdvKYujIR/4gOSt3BS
bAy9cKQ4pUvG2KynoFLxvkB7X4qAI9lob8rQRFhLhnle5zaueHzfNqHxY8XaCH0Lb+GsIFfaYNUZ
fwZ71Wu/uS+SJ4ZBNSY8pnBu1MeWLrySOpqQ7RQZjzKXMr2SQwLqr1FR3WPhW6HtdO1XwOlLmb9a
WeQtz9cAXG0BqU2XMAVNuTHXA8gqhrkpEa4lwYuk0K/IuxOUyAq+/eu+HoMdkvK3OSlaLGJ1vp+S
aUzhUWWBxrRII+khhllz+60iFDZSw6c4EoKg2pFkKjQooSUS76ZFWOOKJVTVMigSc5a0c/jWopTb
iqs05H18tYvtnu/N0Ai/0mmFFClGRJSqksSD7e1ng+kJ3uyejLJux7kdwUG/gr48pvv9qjocHnBg
MNRQEd+kvbvt9zZQuBjkQ6wr5Sb+j7uBx55qB3v+Ldd25gCHvtxsf26yg+Icfw4s2X7KYP1Hf80R
vrjV6XRnkO4jDhnmTmRJVpsoxVyXecLFSef1E0VeXXfscnzYNBVxA1falJ68PM1J4t8LW2uYxlsh
R+fntAkvU8hGrh2NWwxhhrmaE9Xw9gqH/vpINaRRSuOTfHYqDZBt1/eO8u5io/qV4DaoZy9MAVgU
qr3WA6LFFQ8fzEBcaI5bMVrGDCxkr0s7oSrMb0b5HDlQ+YBtrIn/joFd1Y9sywQSV/N8BJ7xPqnN
Ez71LlwIAumDRoRGy7jNTx4EBE+N17ey09rqXfSjtNeyWBIWUiGDYIc7ewN+UtNWTEFZqcSNcKi+
SpZv4F1NiIVwFLWtyY7EJRNPpoMi0iYyu0EBjtURhYkPFU/qg8tP8XgwifzmDXPcrz67O2oGztxU
prIzbaCVOt0U3/4K8hA+33wFpwqY1uc9lFOARpkxLjCMR0jo7XLof51fJp1+GxLElP3dLWzbIHue
Pym/dVvTomgZkjCTdF0om11vHnjUIjqHlOrXGS0TmXa7GQoDZpGFnTTnKTpCKFT7mi2JG15GM8y1
bUm6txE+SgSdPKIzskNWDtBbBld8TPMNXu+l37A3Fls+4gtvBhI4+BFx9A4fHuGofvoAimnMUDt4
dpCTqxk3DpSVQfwH20wk03xGR25e9WxCOxCoRAvU7rw7CMsqAJUcv0SQVOsTWL/I5aCqSHesgs1K
8I2WXKZIs5q+W10kWHXHRZcOnuKJdaoj+5ejnDYyHFhBo4spPWIzF3rt0ZbSLrgtChVDXFgsOpGQ
qqfT212SpeFQzmwraPH3gEoawt6z3iaylvChIihaOyXuDnRcWxr4wVwBusle61nQOOkaWXP3m2kC
7oMrNxryay33oS4UkyKq8fohOQHvP2PkdrF5q1CI0vi2CaK0qXeRvfSdLTkTgsMOFQl0pI3fJ011
Yc3UIH3RcNQojlNbOJfNHYp0ipv7BDL7B/PgzuJ8NwbDWhaR5fNNWlPAjNN2ThjrvvWA9iHyZ02F
/5w6TOGvYHL/jr/qLUfxSgeYZEsaBVZapDmQ+PvrAJC9egavWYA1RIptUOhhokTCPg4WefimFWTV
k6fdAHsxN02+dFYdRwDSChGO4q1Q2J2crbYMw+Bemj15ifa7GHERCfObLhBd84b+Dhdlnm+al0pu
7cU7OtaUSZUyjjBji2I9W/r8YDP0UHNRz22zH+Xpd21Xnh9GkCoO1YlW5Oq7kKYY8OqZ06R6zKT4
QlE2PMf31nU7IR32h2GzUGNQjhybEBQYE3FrRR8lkcZFZ4u3DzzAD3pELSFkS0G76L18QoBP4f+c
efRir6s3U4rhZBi9aYqF90Z1i8I/YCCfWODmfoA2X/hTZG7MmwVbAUSwoAC3bSKMBMlHpMGh/3zp
R2EPZg1CIoOXs/WRE1OHMld4m2L1w3ppqsvKZJHL5cScaW9NSSMXjPce5NRTkNv1SfnUg4mO6lQ5
/gbMRve45EzT9dDDcqIjxpN4D7esclWSeQRV+K21tGsYhFuWyruyVSiKaFMKi2UUlMv+aljjS3XD
RJPUZcB6JCp+qNfdl7YZCLN6kCwtfk9SFwLc1mwZGdJf3Pu4+j4wz4g8R/amj6k6irAh89QJ/ikW
UUN3g0OnNTrpVtDkyaKYlXHLCWmgxR41RUVyrIl7EJTQc+cr00dZPb/d+5HOxxZvbmn9DoH9WHYr
Jv9W6rq/GDVjy6zdxV1F76gd56cKmLG6kR9ThItq0kbVe3VX1ODhLN6nWBiHD3Mli/YAvFzhTXLT
CR8OziJ6EggYRws3cQls4lkRKRjLMiwMe26Cgfccn0+d0LfZe4Jv1nYkQSpIL7chA86YfR2zoBvD
vCFteoMrRFPkl9M33MLU/dycGkHguE/ecy3O2Jm3aUVRaW8l+B3xHR3Xi24awT8IfNZFcALPhe6r
vh9H4MfWnqSn9YFN+jlJ5KDK33yqQ8bNKc3yOdYSTP66f5T6gHSisAgsT7R8vkrPtlz57I2GW/UO
tv+sfwlts6jEWHckX5jxb4UBS8L2kPl5tUSHJzE0TVQLtIyMS4APbI2kc7vEdlPBxxwLX1twG243
UbGnRQjEitb99RrN+tVMdHUuFzsURXVpnwWLfYaeVbs8+d5yjq0jdOmBNw/SH4HzwiS3J+4wS2Ij
AK+nIkzJ8Lg9wwTPgt8cWKJAHCF5py3tQ3oMHGnIPO5cfzwmLEDr3eKqAyecHoa6uJ/w8k5GiEES
itRqRhVVpqheY5kR8Pt0B4BWPJwdxurxofLtuP+EbDXlLaI2X9+R6mNdQKa/Fp2cgEPgJtgcDYpU
DpnwsIkuOmxeOg/tkCn38FPs6Y/QzQa7iWrQ7BgUIxtW85+K/alt0AeJ373+QaPRB1guBENDp/Mu
QjwnC7R5vYYMgdIx9mKyLQ7I7aXv8BJqTDZBpccDc6uhqNGxwlcv488fsuTLPE0HI4PMGTLkiHOy
CGXeSnbumdqAQC5b1jFjiTPKIM96JYHYZOe1ti0CmK2aY7KarSH4RaWSJSCebtV1Hkl3sfTsQjKn
lhVFiHnF42CZDy3QoQTa5e6hOfFSF27DFdX0ihqRSXgE1GxXlFGNEcf1JDMustss6qBWzLklAxtw
QVWJ6sghC5QC77mr+sMNyeto37IQSEkWiCEwCuJ19ycctj5oGFtJ+pkRYEDALyMwM8TF9O7FLDlO
Nn3O18i/gPFgXZiOvoHuUMf6fdhBsEQgkF7pKMe6jYbs8E4NuC+KwIlzHEMhzKs7Rtt7g4kbTgK4
id5d3mOV2ofEYdAEN2/C2ecqpmO0zHA1w3nN3B+ZusyAvYR5G3TqOEdjna0dK/8h04tRfFWYtLTi
vfAivbptWhLiQkFfK6Qmdwk6V/ZZeYamVJ2GhN/QcMPFsqB12uoGc+WrV0UaSXH5uG0CMvFwZUhM
J9lv/6Fqbd5GtswDUurQT14G7UcmptCQZuINHydd1RLrzGHUE7R7u7p1UR+tBn4VYQNHmM7QcqFt
w4F2sy7/XsnPn0RaOKCkAevyNNkVpuuXgc+6OMSdOn65vD/+JA2FGHv8qyjzjeMpwaYgq1kimjUZ
YkpjxAlt+n6/bWJ5/OQW3aQlnpjNCaGe6g7+Etofs29aqT2CWuLFIjVq/bWEBNKYCtHOKJy9K/Wu
6FbbBYBQONr5BjXM6w9oMeXBpFbeakQje3wxF4i6dJ2YUwkNHfaOGjn2mSDKUNvzpGxcxjWcgav5
FZSy2I9zg2iQZaQyVxTNAZW1gZWPJu7DN0lizDMpO2CjpHhjcS/6oSi5I6jBToop/OtOqMp7AlgN
C2IWTkWIv8XUJReWPFOkLwukFa7SYh4h/cQ8f84DzEzUuHUaMC1hNAUi8fUtvj0WG6OlMxhion31
SHNDn0k7BeNrIK3GKKLSK72d3OdVKtUQTEg11cEBM9CjXdJS0OHZBkzNACGaDAuJ4eRh0ekla+hn
GQY9jY2ipJyxQAeQvTwCvHUHO9YmRrkuBNNX18P2512YCPgp9v4Hx0y8bt6kKOUKgvjQA14Y5Tg2
cztfc03ZJsIfhCMYNF9y5LPmi+VcUeIH2EIr79bxu216XdvVyMu/OYdnPtf1gWBNxqseG+GmrsJ5
OybkKtlUQWDA5oOGcOBrBF7Q76amglfZkMJ4150yrWYzEg6poLPomRcOYqw8gXlWZmaTNa7lqi5s
XQAbRadS2U6KyQe0NgErJTFzv7QjiYjZ58UotPkt+acqyLSoTxlxrpLnFMVXXK61uIctp4WkqFsB
7Q2DYsVfxmPa4pWkfxTTVZNBYhFXpPUEpVJaOcmgXp3Zan04jOhiNETfKmtLofinuK/gX92wjlGA
ai8r7gDtxQeE1CyV4tz//Ho69eQsGFVJQo7NWfg0CyeqKLolXVLnqvqbjboRVKVF9aG352EfdE7B
yk7rum6i+UOU/jf4raBjUWcwOHYLSjbUAA2joG6MuCNTx7VF6wFSewJrkGFkI7IeaRKHxmUqfr3f
LPC/eCPg+HoisTSCuezBuIv2PFfasq5TNbs0u8gwdD1fxDS/138zorVi/GniFfjEQyn/c3IKdTc4
hW//bcWSJ8xsCUHMZcgjekghYOszl/QU/t5wrrRoTlCdBDd7CQe94OkpPufZZ3uvEGhBtmfhRgSr
8GdVi61PPXmur5UUlmuDrCx0/ARyk0aXzAVlAVII/O628fqF1OUwMcvPY2GSIj1uwkvA9lE+BYvu
CdV6wrqAX+Ilb5QnABAeThKC0Qkn5lBwWQY7ixWovBTu1CbYQ3YRSUDS+CiuYzU0mJLJcPi7eBmD
3QP6OKXuQT9vIXJY6KVtnWsA+SIvklkwi1HPo2FOWKBQgsdVtAn4hGBEnBRs2Cl0NIzB8dHdqW5C
J48e0k/WKVygfl74o/SKtOCudRLCiPVeHyU+TRF87m8VEu741GMrlLgDQ/4EECp+OPHeJRA6/Avx
74kOYwWCHJ60t6w+U694SZ5jK5mnpOaekXeK5eqzGzJ40/bf8e18P8g1EpKHOlx/IiLb/s3oCnYb
kOjJM+Z1JDVGk6yelBXMsS+++nzKAPZv/InqzxnLTuhYxZJgGjHe0o5MnCfjzzO2waFdHVtiwAaY
Q3U3dXgEOlWXYLbUiazRCLI4NV+1BxELngYXR/kacJ4TQ/vFBrN8qBTNyfq9jwIE8bA323Py4v/B
uk4nYJNWhAJG06FD9W87kNpuZX5a9vo1SHpN/A2Vo5rxhAEQ7zrgcAOGPLFZGZOd29fvt/TE41pP
WeqBRXWqOugrevRT8ojTHyD2W0ti99Crw6rkn1pLQwoIMf0m8vEUyV8bV6JspQrrYZGj1DChUjek
MmHbY8EVw02EawPQBomNYQfB2zrUC4fX/Ekln0yNIxJ48Rwkvg3T6XwGxq4Xl/Ryu9GG9N8Yv+mi
oDUZMLw2gsg37Gml4IxJM/eoZuMzAlZ2B1EPoKANiRW9HSNVuRnbuR5ATMA/lStHuLYq0U1/HKf/
0cmv4t5sLbzSCoShamY6fDEclPH88D2W8S1TXp+U6jqSxPpkYhiV7duGLqj4Ys1+NZAlh3xTgZNK
AtghITzUbJtVLrPBPDxjtI0wlwa5Ns0dBcS3Fc99IILlOh/LAaA+CvFPo5owju1mLBXmFJ0qw2Tx
RkCvDemAaYjHNa5ByC+lJLXnbdj7S0pF7ZhUdz+LBSZ41XlWBSjlHmHEFvIXmz7XjztPV8LQX7jA
o7IVQw88LoNy0AB170wYCgh+CiFeiNqKEpBiF7avjJwY+Xy0CGW3RoaqAy4ugaSaeTcFsKlV0L34
KfvNDZcqPyqvMITLzfkWVVoBsJrj6TJMm6883/vQ0EiBbTM+OGqmCrMHTvVdYY6bd+kjOBp2isnJ
ILL4FDHEzzYgICH6nkrgfl/iWgugUNnhs08bhJvK6FY0jOKjHxPUPQT6aJKFh30K5S+j78lQ7v7r
dXWJbIBSkCRga1Z9m0rfNAZXGrzl67i0FxtnrMJDDaS19UkbdmNXiuxASFgkR1ztrpkclM9fgEwr
rdEql8Bs8n1AVAAIwZbeOktylIkRYdbIgj2peI/bUsmf9H5yCn82DIJDInEv2QLTMev1PgcSzc73
bBhNGHu6JGpCY5LMzUeWeluurLgGYdMYubTNCQwhqPO6CjEOJghvJKb4g/BBwC94dBN/z85Vr9j3
WQ4mY/jIdrZ1lVNIrDpk7iFrVbGfez3MWu7hCql0oalssu1CZG8kZlBa/Mb9j0D9dTlQ+fVI4SBz
sJ/41x1uPqP9ZcyIbAkCXCvChAjgs7kLZpomrt/3rC96Vec4yg7RgOJISYkLdj7rBuiRq5p+LTcu
88eVnHgEB8q52f2Xanp5LedE6mm6g7OxXqiLu3erO+K55SThRKYeBmcYQhBolKLxM+Xsx0haNVN4
wNOTa5S4z0R7u+1MGiRpwAYHwN2GO48JF9f63AFFvf1hOElWANpaWWya/IR0PB+4OOPbG3gBHegH
V4El0X/T+NyWEEDvCY6EYIlV9UK5KLe6jp/Ye5qHMtfqQNvDx5D469Nf5sMdGgwLiyS8Ynd56NkA
CvKDo7lp9Ug6yMpfIoLaW8tkaPTEIN/MTKgsSAWu+VN9kzh/VMJdVbMJclSoWUGxghYhmUe1tluH
dt6Gyds/ZHmZItaFUjaHhq3PljSf5fxQNb35MWJp5zwmkRGUC1Yv1Fi7TFt39ReehcBn+Xm08T3m
Cid7swuC340+dZXqA0eqvl7dNCt/dwrU1nFm21gewIHis37lx01XxHyuTC/rF4R7eIqfy15UUWq7
FhrnIPR3JLz//SsSOclhuSUHKl4UUBrehvzrFlQUi6WllxvPP7LvD3EReTRwtn2JQ+qWtRg1hiqb
cHUTc0t/Bfs5bnU0xFYcmHBYXFCxyVOGo+W1Q/gQkCcGjCczMDhBGUn8Cdyjkopfgq9/MsaDezqM
E4VF/xr5XtL25R+i1eDc5y/KB/JUV44AX7ikkzf4kYTGKu6/e4TZhKi/rt4+nsIFaU2wvkERZvK0
lBym2AZn0+DXXlOeN4zKoUQJWmxMmCTs5VtjRn0VM5bHcGeCGkVgrOMgAr3U+kKHQA9d0mZmEtS7
N0LoKUHE4llR69sFjkfLAvzkXOFzIH64CIBIXvuwE8OE6GsM1FoNsubd1zBRtLec24ri57shz3kF
j3Xs/CbDl8xkSucDAooWNl5YyJIOfA4v08G77i7wiE2PzOrwBE3Tz27J33o9eIZHw/1I9mtUYXFx
xH7dHZ6/eTWhgoWjKC4gC672YQjC+JujVI5q71BT9Iohm6RQnjijqy9/DcGr6hsevtiLq5MtBCMP
U3Sr9z6RCzX26pjqCNFWMDZa8kVjR0qRXCsPTYfLnw0R57Rw8vuBn1hBTvHHuulro2dUOGzmZSNM
7Ow9TfpN0vwDS801CGLHnNKwfyvZyD4SFzdjpkvont0zYnFliuoLCYc3fTu6oqsKDhOzZcqi9lwo
WGIeascwMdW+F0abaq5OqlPSAAqRjUWMYV6ONlMetaudqSv37LrWSjvdGilNv25HIvWAvBPrdYvr
aZniLIbdBQdicYuH64Y7iZAsnNMNW9eh7fXJAYSSgpvJqH4lWvWCzLr91u7DgH70U28mYyEl8L2+
rh2+2x5lSyPgP66wnwV1TAXGYhcbjBuEADGo6G+z7A402DdTs1Tk/PPSE1wbixThDnhHhid1b4/q
jxqTFucbxXOMB/DF2HGrVKPYMEWln+oR9awOjoXUvg0PyyG+UcRWDdxQWMownq8yhjWdy3ZBSGev
ioRhTqCP6SQCAP/x99ReQ5xy8EeFxUQ/Dd/fJcgg3aI1ru/mxGaGn+IjJd4xyaMzPS8yNeIzyXSN
H1CvWtzXZYZlOW0H3mAEigS0YgFvIgTq06naFylxrcE4wyMBxzWszZAM21Cn2RSe2oGNUE1ZjCRj
UoBAeoff02JfAfZ1F2KzMETM9XIjizbBQzfrFPerIXyAfGgcrFH91eK2WTSolTqyudAxrDDBa9vq
ik/qgBxDvd370o1InQCvGfA+Pd9GtDIO5KKKNzGtfelL4Ot+tyco8TYO1qLIW6kejWKcPY3mAtfA
d8E9yvLOgenYFUVorzZY0IdDyLJ04dcmVfOSjFe2UiWvVudOvupezWE6h+0t37pz3OYsAEGk9eZM
3XwBFeA4Ypo4LpsAVBKOSJd+/s5GsRQVJyZWg3zfQnnlz77ugG1aPFaTkNFMHRf2HwV2qXEDHgzk
/jpCw/KFAJikk5yGdPOE5jSSme4qAb13v/gUViNkXWTg0SB9THytgoO8us1lvzRWtT/asRDQBwyW
vA07lhQvx7rkhFpq2YeDRrFtkeonAKAPqkNkGIzSQ4xaLSON3Z6X1UOhGNEmgx9Hzlu3WEFPeo8b
PzF3KuiEl9h9Ej3XmPa/tVr6kwy/Bt1RBtSgnZOTe9cPY2P/KT088bd3Th931qHpTm7OPIcgT3uO
hNZUHGo8UJph9/CdMCYDjbWAEcifQRGPT+lxGQualhTXVJFJc4MV2n1PlihvabWWWqX7m9iWP6Gw
b4nFX7G2YpC8nUrabGQRzvyZk0FJzLq16Cv2Zu5ZiQV3wyK24I8cJECOC1oCAQgyT15IPi62ualV
Vo3fRVVf7rbAvB0sx7AQPz8NDTWIPbL0OqAyCdLvR3dkgQiU4/gs67Z4my1vlI6aA37FbNKmkaVp
x/nKjsVOamvWpsgkrYmGwUeMUyrf9xD12DDQ0vOET4oiBsk6Qc77/gOdKHgXbzbKUK3SQSkxej9N
czQDmaEfRZNdN5kcAYCzggBLOHsFudANDAMpwlV1e8IAgpV4YXmkiJXUX7lxOD5YX8JMNj33EmlC
yELbDvLpA5RojYeDPeOhrnfkukZoGRczRX2dooyGCGxhHijCA8Q0PGOBS6MBXzrry1pUcDGd6b93
CRlaVRmS/QPeCg3eCBktoBtAhJIPYSD5fDzPz4nWdipPWYBFVBhY8FoYETWaehMrJIX1TBWAODjM
fycQWEK1ZvKmu1c94R1XoikH9yihbfdHNIVAJuK7uVeYpFK6p2ng1vMzGHKL68gWObiv/baQszae
Ud9k8A/5t36G7QUPhWlmMaJ/8fGCSRaOwWCv+15c6mE4n/EmGbSoRkiCYHc8pmLbeQ4VqLOA1oi0
8a3OIN0UmbcVtAcFoss/GMNRUYKI0kQ+eWslITUU7b3smi6mWO8gpqUehQkkdVb8MJx1F/MDd1Xr
CpN92TU5mCi9bZ7pgf7PI8C4qYUZSJfkUyS3WxHEZ5blq3FZFKDtvx0x/evO6fLxi334krTWWtT+
t0r4fCU4lzFCSlVrFgJc4BobPVdZioAlLfwoRjZga97qUsyHVbe3zaIYWjEu1bRyn2KwHj04RCbI
mmgJS4iWOFRROck2/ErsX/s5EzD5GTnQzz3/x4Vzvl5UwNtoxWv2J7Gr7dwMkZlErIDLMAdfS61N
EXqpyL1TrKoBWyowONqV1fSKL+vHA+d8T6KTqx7lgaSZq/E996kIGZy2EGud/9Ir4yLZZTtTwhLS
ly2VdQv6oqo0GO43Gxx1qN7wNBlPeBi53TPXzB4y8J9PhbQYTzPPs7k+s5txSdQGmYqD1S7CsEdg
qEnTn0MsAKQDzHDLGmuEjBgJ6OXg68J3PGDtRjWNyKaBR4ULHOkDptJ13P+/emqHP5ZNKlACY2dz
sVeDC8zUhpq69tMwhipwP12ykHx8CrTrMHeIxyEwq7T71e7+p6W26io3jhSfXu0lhdaa3gKca1/5
b4KwveuS4UqO9oJfHbjjZF10vqyhRi7dZ+9KXFbzaWmdCuk0PMz9r0pV1O9Ja56BpAT2vAZEkDmy
zhgctbrHgmcwyUILzBC0IWdR3fH63AF3Zb4ccdf/RTpvx82djVIc92vitKfbwUZGGRN768kykcui
Y5Mh4KtpGroIYs2ZemUo1Puf143Mv+Sz1SrLRnfrBbiXa9GhClTyGfSfH78m0CNMW08DNd1icH0m
ngm4whto8IcdEf9l8mjzGmKOZVu0eOCpq6cOqPnxNIFzZX4l67VrNK2xF6GNCOXIA+0IPeQnUhvu
qCBIurXxK0qrR6Jrv41FB7mbakY3teGYvkQUSwvyk9quZml6fYx/1v+nxqo5BWkWsHNTa53x6CB7
5QW1ulFiCSBtZHIDXWO7ZAaGy/irb73SU/1TAURaJiNruM2edYW62n7TqmKpww47pQsSdWxGaPd9
mxNHnO+JKrTUDSLfT89dHhVfa8BKL/qajfM/XYiSLPuWKD2Amy6r871r93nyLPI+y4QxLrp1F6gi
i4XOfDkW4M/tU8HNL2DRVZHwfEmWi26FVSyKhIHHoJ5NA5QlpvlCHjMmSq6tKQP6fhdSine2JMrn
9J04UDPahCXXBJ7TRIBT6IAF6VMhKhLtsfs9x1lkG6e6SgIdgQQrHHi4SGGmr5JRbEdaW0L4VucV
J57FTKWX2pMeP1Y8Om8+IoE3cQYwRQ3bdkQiIOuQpEOni8r8jDSeFmsI6yoHvna8FDvLXrdcP05+
28WSW/mEchVqJtCe2/QA7MsYnGAV1fOSfKUG4AdVn0eL+l1LXPacYeYFHc7U0NKkiCs6IAWxF91S
EaGEadRXnDd1j1Iasmogi0l0iBm+mqStEBAou0I20F8Ksx2DYDNv61vSZRJl7Hcv9amr7vgdKUce
NBnpwz3QvOOVqq6ExhKFW0YX1N4eXdOXXUm8bP9D9XISSBh5f4NnurNG27HZIJTtTDvmuAYkxAsu
4wJGpPEqPoQnbfTvjKSrtldHrB9BmPlzI8tG6x590qPuCY82kkxCcjeoaD6sCWN2QmYouKsg8QD1
Z1grmM8bWeF91/YORo6o8i2RIqwIqkUuLY7ndJVYkmKULqi0VAZuPKuqzDBkIocted8Ad2K1RFmM
dVCGmc3+ZacWGgkbeRmzpYRXHhjJHhY17Lmnx/6NnVs5bZbE0HW4b/+2Y+wYEPfKZny3wEUchkwt
Z3IIuZad+dJBSYhM3zT9NhfXU0k4O3US23IvcTPsaUMKjfOqsir+Ke98CFfwNyPFFd9Crr0OCHll
dq85XW5wONIkoWgDav0tUSMAr6HRCtdPqhWT0vT+Tumn6yi4bJ0tZ4bp4QGm1WWMwUuGKRsLLkpd
Pseaa/2QvZcMbMYsCGn+P3ZJ/YpjEl56hJbcPWUhqGu2CvBf9D6UAs9GpmtZ7yZkT6gWvsL/OvZe
/XOblB7qkwQNGHVXxD3Dwo7IlHrT68+RjUvAdZ81cQAUSCsM5NK0xa9kwXeY/utmbb7c3boa37BP
a+Q6TDwdoaIn1pJRPGGiy/eOmb6dQ/jcMOYkNOU4Ws3w0L61y40SoNRCamoKktCK1XXakUGjS7+3
NIhKED+vzp6PORveLwyb3HT56uWMGKMNCA5Q6eoUMep2PAN5PmVnQEyWLEnI83lEBtCY4lQCeJNt
JVYtztxHFIKqQP3X7uC/btjRrMMfQ8f5gnUqLSS/nprHkRAU394AIpSK6vLDkw71wS892d9AONRG
RorO4GH5Q6qdqHOPHgycWN9A9qhIqskdzHWbf1zeJh7vv+E8ld2O1JTYJ8hHnqhOBlTa5ovCtpOR
T39TbWUmficETtMqSiR9umFuU+Cwsjca1i8SugZ8mz2Yh4vCwCbWZZbwSzPcGX/JSXSlJrn8yrzT
kLaCkHWOvOcwwNKBen/ZcL/Yufb19ek0fSzugp6DqFKgSbRMz2OMHsmqysvjRjm13L6HG7snosS1
ke3lba7uc5QRk0WGjmGUcIR+MzlP3UEnFhG3uRXgiWNnqI53JNLCGKotb8ye4epSl8LvOfykGHw0
uzZ3Fl4QEUjiQtup6ONBWPI903cz6rHl1guGzS0MiIBhzWbLmoOU/6LW5Y1hdhn1J1WvNF/vP2Fh
Bx7pTiyY5jgR0E6rGcEpxaaC9EVgKs3VwpPM4I4VPlbmi5soKgiNaz+xp1Ds6ej2OHLGFgIYmah8
IodBPzorPSyqR9vOvFXKOuacNIs/3JTGhYM8R8Glt8VTbw1yG06KJp1tzGfozw7+aQ17r25ap4rZ
zgl8DvwGwH5BjPL2RkOASSeeHL0EUWWeDKMnrYwdTGNErDYBe+Zy6VcM8+aY9ITUmSVgHDBaHOZU
NN9HtgixW5egXohjk5PWej4l4dzPF6+dBw6CR4HKPl4gaTD/aLdb60SipxZp1waICoXLbN8ghwm3
wTMTMWcPH2kKM4QWfV+KdA+Oo5bNZVWcq+EvnpkfFi2WUIbLEpzxAZc3aRxMVoDuJeW5s5TU0sjE
vS8ey4bWdCXxEUVTXANON0kw7T+Ik9TOHa5bYRc5Z0TzFGeil1GeBMTX4+tUt3U1dTsI8rHbvfzw
4cFv43xsgdjrMYZpWtnhto3958jYCy/+8eDVDeDlvVQVSN/lMwMlNpcPygN9qyaExvhQ2m8+X/G3
h8SXaWSkEsWMo5S169UglR26Soq8UyL8Wmy6rEbnZnkhmVrPhVy3XvEg+LfMivhUyo7Gj3OsDkhU
xyAZupqbB7WzCKxla2jvNJdj6HyX0pTHEDOPYFX/vWXWaWy5Zv3XU0vkcgkOjvg08y4hNbrRm4Zc
AOx2O7EFt8NxPIXPQObzzrIXI7/TwoyKHCYLdYYptF6aIpXQTJgK5noM22q9L79e0zGl0lMMMAT7
JOdpqMbetIU1fOMaUVUm6wqLd6rJRHzVu9zItDbku42vKVvT2agJRUvjbKJX8Ixemc7CKSjDi5dg
WkfhGp4faobWa1BDholmpp+Loy9Y3yDq6BfluPhIVVmGEev5YO0feujrP41iyAjU0ccoWdSsRPU7
cwd2YfMn3K2guRbfvvzi+O5fM7hrk2MQTl0lgo3gN6wXTEFIdG+RmwzPI6Igfp0fLbh8A12IAHuR
YGkGapHvftldYqEZA0FekLmthmwAFaGOupWwm8lZ4z0z5Dwe8eV965NJQNRz7gt7jS0GRBv1zg2X
5iS7UEx1iye/QJQPlGfrseu6IPHKhXagB1A/+TAOvfcdinNocL/i5m9J0bNkYjO6z+LaxdHjqygp
OfGqyf06/gxxqSecBEAe8yq8fc6H0IPtlwem79WrfdmA4qOhPauy/x9qBqELUsvEKB6vORcJgFIE
Pyrn24fDG7KMLrdYEyhgiuxgPymGgq1mftn8q9JR35p6brAPMqwLKGI3+W8mnVEUsW6X11QLH2ma
pnIkmGshRwtXV1osGEOqTxIjGJqNbgTXuLHKYAp2vRoElu8pYTP6dLx/tQKDvH/pir1h18hnnv+K
6IRmyqz5njlNYJ1ky6ftYSG73Az/rjFWYXeR+AZbG+zgQQ86MsKTxXjVqQ0T9T/QUZPahngfD5JK
b7d32WQ9AO3MNGe1vDUUWJAzB89zgxINg+8gTm5igP3UQsTnDtijhcsl8GpF4ZyC9Vv0BrAKwfZ2
vS+obst53iMmMxS1Xgssym/iQeAhIOTdSs5fW9NQH1CGC0dO0R4Ng+MN5ARJabsIfBEHARo5Z4i/
hFMfUa7xCzYDXi44GS3OTyl5EuCAMEVpVrZg1JRHOgk7AOgVS+dswl0/oE0WpGXZiLle0ZSBI1RO
5egZIgmWutvGwt193nfzw0Oen9ssjJTlD44ratpxQAixQxuJao1F254lhLziwG2Y+yf0s3GpadDQ
stLj8pG8UB0zT98i2E9k18t0TQCZBMOJ9w/3vORqsLGfMlVvgUKxn0O+K5w/C/BR5JXPFhgJyMD/
1ohBGjcgDkJ7I1MREAnYOMDWuS8fqYZ+JuavPmVSvj1zb7EGy4uIFcwdhqmRBbyDJ8S2Z/qvQD12
HOZ6H5d/wkP7ss8ajOIiQmi8OLP49TMGXxjwirpllcFEn6tCVeNEysgSlRXlMnlz7gEi2XwQceg4
3NeNRKNfndgbkjelB8QKOezTc72P+hwL3UQGQSv/O+U1JcOeZXg85h3CXjI30pYvTlUH4kawDl42
/mzfXjjEJ7oFl8vQhGepuhrmpQpA9pWowv/YvagfrKCSlJaiyOypjXa04M9FnWn/GjxDU4E/wcbT
Wo5gQgiL2kN7b0ZCak+fqyodnbuNWNPa57C/aQMKFreePDgc8UplLew2Z2r10z3Lw87Obm2g8Bai
DHLY81rUBNJL2rzivvKjEHM326EYCdh2v1dGkZIG3iTvogG95nmNhVt45iAFi7V4sZMz17Wz5O7y
Uk5ozsFFN0Ke7VcI3cfLjnZfG5/wqcgR7cj7CXk/TKd1l998ESG5Vcft9mhV+TgdGXI6tem5+1pg
LLgraG28s+/qVjZIAfqU03yuMtsKNl5MNkpvMUf83MlADgbeZCPuhB8nfkM/5AwJ67cjOfrzliJO
yQ8FDzPW1iou/N6rSN0g5nhVhebt/bzX9wPTIza9+i3ijsFzFlDsHE+RH1nfRXG07XcljknpgMEL
SxzqPdmmeT12oL96L70FsNxwjkn/GGpq5Mrq7dZOZdEryzmwxth+HbO6QBe/kFRAhdqlbWsH3sP1
rZ/O+g9ZUAxn/VjRKnXkP0eb3pcV6IhAF0ZA19+xOn9fP5s9xNCzzukkMckLnKa1EuvNBzH7+chX
ZGlQg1DEgVtT0Xo1YItWoUxGkda8s6vGw+Io3yAjG1yv0fTwFMAEC1CRdtGJYTNIU+/U1m3IT5oi
OmcH+IzBUaof8KbKYcyEmP+ID1QSa/45FkWQ+gbspKVDUVvhMC6YjiYjimPsM8cMGxcqmCgU99tc
bNHFK+LGRD5MOW5xisbC0zOY+9ztnEeMH15Dn7isni795w6yZf5/vMAXReDrOflqOvlJsBvGwB08
Bf8GkdCH7OvSXz4r0w9gWv5pTVgnp0s9g414WkmaUBD7Fe9jmtTl8ztb2KdtTAQaifYhGB/z9E8S
aGbavBrx8IWlxRWXlYZNtYwZ8kAlkYKrrXwpeDiLhFRcuHKnUkY7uX5Hxr+kf7w0KKA3eFpcF5Np
xNjXS9emHHgsFIYlcvo7RWNiftxqLZMTifSIlG++evjHuTQ30dJRsnnixXFukhdquaw03e5QIW0V
r9JZwaVdWtCQtTEYrDvWmljJwP25Be5LyfdRkAWZwfKud6Ns8MyQJu+uI56PFgaVdVC+FgM+Uve0
leAf38cn7ifLOZbbacTITAn8pdpLZq4A/ZqL0j/CQAgHRvH/MSGZCwgo3zanjHfN96b58mM5SNhu
rQZ56+hMy53pPS0hlL5S7qdNGByeJ43jOu8BB5OSmlfXg/fwpmBw5v98B/X2yGvTAub0kGCdatLo
4WkQz2Q+0DdE/yJzjvIta7/nodP1ac/jd4SphDjCmRNVvDRjh/biX004XBgFFAR1EDZF7HP0fSIF
EfxAwGZzqNTi8FJRKijnW53PafAmvrOvJvNYKdaMST5z7Dt8b4xGZNqbqWgXTuNpaA8sDefyBVY9
TbQ36XN2WC7hfF4njz3/ms+oA8jtMoxMuqbKVfyZH7cRPfskvNJ7wyq9IN6Uec/Poe9crSbQwKLa
TcRIJni4PhYmffJCWie89XpBLFZcHes0YG6xQ/xgOvWl920KsRNAkcGSmljTH2F1ZPZKEXbLeIPg
a4xxZ2JWfmVl8Un3BIm08LyuKIhFzWfC9OPY6stHeq4Ljsy3gZB11wEk7/6/6/ny+KVJw6Omeszg
v7vN71Tj5ht5Wjl8bEWRd87Dne6xwLB2OLwmBHFdReyFkl291mboyQF0Lr6Lr2qMCuiW58wofMiZ
GedIRQy2WXljPxAYdXbIRhneEfSOWHSpkjhu9jf4wc3UAbZu1twVQ/7XP+ixVjAU2g/gVWhy6dwE
m6hUUwvolcaxGwCmGr5MFIStpOgI4WyTxTPvw9IdXVu8W5I7/OfWWmbWiE1JN4P+tl3GHlb/pKbU
Hm8cd+qW+vHdQIbu/sSAS26n+Wjv/cDamnNwK1ho6vC/8ucaNNPt+z9YJtJvzB2AWqBO2dAmtSo9
KiGY5tmxpQCQ6X/B/ycHgexU5k3k6nF7ZMkmiijAzcXSGyXvFjZtl5/orxduIx7UaGnbws872kSM
9SVlb/uhB9vr1gGu+kubuMzhnsu3+qnRXUBHq9j1Vy3TihzTqocKqPLJ40aB9Ey5Yccj1nQAP5AK
JVfMxnwx4SO+B5BCssrXQl0TdwXIdu1xBm+39WCYtD9GYbnudZ8DttL97x+CTDZTnwar0s8wPGM/
DjLmcN6sTX8dFkvfEdTirxY6O2inRzQrp6B9M4SS2FFUrW5ryQZVzINc3bksZnHORAmHlsHJ9CLj
iRRudxJ6kfWptOXFhQuK/o93xckv1mudmmzH8M+xsUtLiAhmFreNyq3Tt1DVa8rwlG1bEwyWd853
Bz7l94Ff8jNHXJ0gRB9TPfLXPjjRqIIx5MRpCqt3lO2217b9i7HlJXa725K7JhHxUt42cwLPsJZF
8jd0+kpqzxs6FJm4ayjNw01EqCbsDDCwrQhd1od/Ec8QiILvhoWBOi5C+AL8aMaZ49yQUbVYuwTF
Vuw8kBPNgjAGRLVB+98X6S1GzO98wNMVhAdYqiWHFDjAldG82MCSt93+AG3/m2lOHN6Iy8Dj7/o3
cIUthKgbvR78e7ENLoLZcEhc6DjFPtcDRMMPGVat5adw7Naw8xjD+/vxI/3rLzUAWwH7O0TOhLNK
eqY79tYMqQQCjP2qKIulvQ4WpTjGt5DKYXrjFwmdHg6+5k4If8fWmoDFqjtvB9MrGyPua+vM/GmC
zgyVo3Yg6Ufb7qlUOtqXD55kJP7iljHv/pUIgFGZyDup4HXDQ3jicevfcQdGqzd/Wm8YPIBMSHWO
ENRVhJzg+XVOqnpI8FrF8rCCP++ZxaGk6JEcd8iZaKZYgBbr5xo1Nvxu0U3tQYO9aGvvwQoAjTJH
Omy0jMMl/DrrjyViAVT25LXV43a4Ew3Lr0Xooa6ORmNkeo9dyeKpd/OJjDvetmZKUdUfLLAwW8Hz
uzwI9e+YoMA5f3PcXKy1NXi/dg9s5GAbwRDavhYNTJFEn5IfX2jH6qlupdSEtXCdx3JhnVkYHbRl
+3Vtq+KGpKfixmyjrBaI6XhPnap4FkcBYX1O9z9sN3BINg1yn4Vh2b0fRoQ47xirvhIxoPnSAsOY
6Iyj5eV/rEqGd9ZlA/1xMTQjBFhztxPzA1GFBYHRM39DVZQ6jUsYAULFKVS1fhovaDPPjxjZ0njQ
i0mBrCJ3UxEFQYf4Ue4yV5LwkKjU8nfMTQ1ZP1Yx4gA2RtdCSXebTi0Q+ugju4Huurf0BAktm8On
yvAvvrb2sNXX/N/dR99DssoElUoed5/pjcw6zocJvrpj4oKmSJFOVD6AvfdznMTVAAwKHqarY26l
jQZB4Z7q7USimhxz6TFD5QggdFrz1fh5eTgl+1WeOJUI31ikzLEJ3b8AIHXtwSMhTEjbRpsf5sCF
UM3mI6HqM5cKf2IrNU1e4XsNpT1SMNrvHQ554bq5reKaWHqcBi/05nkhGnwercv4Hy0RKNbCfoCk
dbP8WrlBFRKvDQ/aA2f2VK+9CbbKEbexGAkoCcMGv75ei08ab8xGZotI41rm5rhRJhCSCCAMixYI
WeZcvQgVKE4Dmk6CaEF1vvZboJrViR6OJdAgeK4jR4ablbgr//Fqs08T5aZs6LI8c2UFnxDOshyj
O80jh744OjChFAJUlpARABzB2krJNlCUsX2++Vb/689Oi1Jbd/z6gQvPtfdLUnt01oQ1GQwD6HFI
Md0rtMzQLewGREscdncbyJRxtv1zH7JAe6QQJaBMiDcYqGGhyH5456RdLnfAMV0hh0p2X3td+9mZ
vj96RHhV96ypGtDie5oK/uEk48NS+DNYO2YtxzPI5Kpn3b3aomT8Gbl6d73jHyYEIMyvLTfqbe7T
e5rgK4zKLSOHaUZykh92cPY4hfmYvb+U42bJ1yLgEkK8KSszBNxA14F4ZTGGSi09f65muvI8K48C
5PjFAxwXWOTiIgBSIXCArXI9QTUCK8a9fx3tNS0st+F11eKA6Wl76qkrmEHmEUVw9ZocIn/iMQRD
zRjqRcvRQjeBfkxc1DwgV9Tfd0e7hWRlrPzWg83h1m5wdMAENnwkoLJc5KL82BaqFSbEyFH1dFlY
P0nnH+sb6pg89QGIcuDc9F3b968y+BCZivtCSQ+sP6yjOw1OporQMKgj2nEcPZ8dGLUm3gb+28oD
25aZLlkBCYNM2oWX+PxXPYU0bdnZoHZjpGMIwVQgTWdZnPtlyvZqxNz8O1T+yU8pi5jJpq5/4UEX
Flqd0/5BezoFG7QXzyE0e0twKOOnTtae+wDUzN8BrS6KlLnYvpTSFQ8p2DXNR1UE5x69kSiY8XdW
wDAmCqXZa+z7PSt3od1EYsrjPUeLQ0hT7WsmgEG7kDCFZoMbpiH9Uf+m1Xpc0g/6a3yfrW4jX+eo
QkRdl3Kf04oz/NrqYcaJLUhEGF4yJBnxcPBEmYltAmY6cHXSu2tCJWD1mknIozQdCSvNeFZBsxNi
jfb0dEbx938FPjEuYGq8vo7qAhSXKX3ek4xj4FUFNWzJfF9N+SrS9Jw+O3kNFXdbgGJa6xcZVokr
o0E1VUAx5RDFzawGwnmMXrSQBaPO4VpCEvColMe+2QtuZ0T/Z7YaLR4ICCwyBqwsfLDtNGG9ySJd
6Bet710LIw19/iqLc91jb+kZJM1w/yQQncagowWba3cXw49n5O5NcHJolsryNuuTILypZQgvc4xF
JGuXE+PGWzydiMDpUuJf8CId2XIyRG1eAJknnGDOYWr50y2kK7e2ZQ1aeI6oJNslYQdlT/TZOVSw
GW1itH+6k0uOQHgrrqj2fRAmlmYR8WzodxW+Rpy83kkkJEiomvDdddw7LQBwJjXMJnwCS4vZFdZF
Q7jfrwvM4Qzh9TzRHT0pcM2z7nZtOWslBXYaq1nUGn/xuMHkcG1AI9jBik4W9kMko1f6ShOQv5s+
loVeJ9VIfUYQF8SDh5iAf5hjruV4kStJxCk20kbeoffkEA/edsNYVxgxhKNIXMtgJZ97dwSL3i3S
v6H9WvRUKMu1OV8CxXSwwXjRDfHJOosG7z4YhcgxY/jP0gT4QK03IWdGf4xevu/5jqQNhy1Z4aSO
7flj29XONAD+wN2iyKIFmUUG0VmeTm3ewcidWyAkqmZ8Z+ujyd38wQJVlAzkdP+Xo8Q5vB25K9sW
bSVLC/sVXDEXgFUObymKm7d8BZobAQUA/5VTsQbTF4ObeEv62dHKJAkXaSb9lBT9HgvRIl50fmxY
QVT+d/W8e3Anu5Rx8rsEFs1mfa6T0L1j25P6eXb0kTJzyuBNHRD+RsLSJgA9TtaHLocxMr640b+p
4+VGJqO6/ZzNVC89mZjd6aFMz3gZ5u+85hxS10fyawDOmAKrjQolb9ZzCsXo8Q+TJckZ/16E3KEb
qmcxxDBgSgT3dKfIBTUxozD1cF1tvJ117tzqAD5/so0LckRu0Wx0GKZSRtmaDCVFDPWW84RakqwX
9BGLwu/9ZmDCyrEzHLoIX4KSV2uJiesgRA52jbRXUIMJpJ7zeCx5qoKoGEhN5qPSAy7cPH7h6IFV
F54SNCVLMrRp/0qCm6/EBzFX+Z774MBHoq9Kv2Buys4zZnkHB3IuQU9Y3xzWNJjYYtsjEEm7AYag
9obiDrTyEecBbXlIYBRuDClsUxP7ySli6JUEpGHIjj9VaOj/KPJCwswBWYZhqZvCl06zDccWPkWB
7qBCY+ucDr+PG35A/qmOSNyZ8hYFk/C1pX1y5Xq0GWvStKjA04ty+W+DZWbaSrSyceTzd0gAXtMo
sWsG1mg284gfpgNn+1MdwNxqVsub7Xb9+T99MxonxHGLhw/XjguMuXOTShsEH0jQCbBakcOalajQ
tjzm9qw0K1UQfWCQ7ctUtFHjeX9J9IU008oXI1eHOeNA3ogR9v+SuXdoRMm/8b0OHb/BKglU76yg
c6A8XMlQUzXsM727/SX5MecWjhUCYpixxDc+WCYiU23a3NQr7GsHw5HXx88t+SwVbIg6mGBaYaWN
T0qyFWwwV/tNe07Zn9Nj45ZdmSUodIgdyWWik5gSVdr88J90wZ0M1Ckqe2MDpx796+9rzYPiJM8G
0QTXHU0Vyeg3Pxiyx27QIlOV5yCDKzeOf6xC6mvf6jqUK+Xf9CTHmc/qJ78JUIXgIS8w8APnPL6t
G+XdSYG7IizbzP4OWcAa5DMO9Z4+ej8SpBr9p0hoau4y2TT/LM+87agCQ7oz/YNKlbiv/QWEKEtF
JoFK6qvpM9qJwfl+rhD8WjBd2d37B2d2607sOriShfUUSB55NSXxmV71mt4wHTtcRrBD7wVUhIf4
FmEmOPfX3A8hsFKQoVPANwjOOGe5Gt396kGnvq8ir/usuI4i0C+KO/MF5HzfhjYV0tMxlzdzcY2h
4EfhBfx/rJrBB0D8m+Wr7RqJaTbx2PCYC3MEWS5myb7sxPkc2Nv084kz1H+W3GyNJf174/Dxmsjh
44U7fHD2zkog8tq39/olfzIFpCgSgz2DiQ/RiIJ89d0Xa7VJMbGH+1gp0eazsUvwAMRnwhPawEi+
hMVeWFNDWJOenTwSY2OSQP3uL45T7jniEuGjk2kx3aVfTBPHddBmmRApei7fq/qLcICOeiVRCXlC
8iTbjZMJOxxjIXHHba+tQis+YmeZ7u2RE7QbJ7RdynCuEYCey8khuYOirEE1IB2zQWo2WsAg0BZm
LO97rMxMsSEF2aw+o68wT+lYhgWRdgj3vyVZ/QjPXP2f1yCzSdP5BNV0gc28fBYFJrqBqh03A7SX
8QNpMu9X45gMUo8SqVcxkBA6K4+GNY6Hite1lsyV3dARp2G7WQdGMhbr4KZ+7z+CFFznL4aePOy1
wQud49zL+2pDT5ohlGWLhdHMOeLkf/O9NlJeK78+5L7g9gk44RjDhGBWpYPABNMLmeqmXW006QVz
q0zlKnB0AM181FPtlKJdoqge0D1WKRp4FF7KQB2S2EG21+ZjzjnBrFsqjKrA+oFSnJ7xJIF1/Xdb
GaoCZ1iwtiI3PeF98F5tPlaJgt0tzcNgJ8XFDPZOXkmozKoqshRYdmDOD022D6GfuVRsJ+9w17R/
ZA3DoSgWVkUej+Bm32yfmRCS+W/CZr8kY9aX+rRazLRAgNH0ySpFX305B0sozPL3t4BOCdjjDUDy
rZYYV9QUmAWE0yoit4mDS6GQ51tEKFqZ9Iirm63EUOBb8WjB3o2eFjgRLVy2g5DpfiPFf0a1UEl7
eiJ5Ks1pthrg+qukms7fsitq7Gc/8zAjt1Jor0dSBGRyFfnTQNPTdxb/MC1D+ifhu0uXEH0yl66z
9OoRO+qWxmnGYxAAVwB7rij2Za8qSDUUETOkIx8DgUaeLn0ryyg7ftrCO3Udnp52BfAhnlgkFcgj
5akS76Ab7ye0KVv2p+/9yJ3u/5OUSmExrHsl0Of6HnMvYDgZwZo1ZEhdq2K4ks+j/F0Gjcnmwind
DAB1ijS8AXITmc9vEdYBRnydT46Jm1V5anhxTFqOryeDDnBsUXZJULXjIaZS2iLqFthcQBfqRdLR
Ik4IQ9RnUFpkyHAsWwahLUJ5jAhSekQB+vzGoX8d3Ag1T14FgaAUlFRr3Rp+UhK2WKnkQ0miYntg
Za0Hse4/zQxdsizWUnJ92WXuQ0hPQZjlVFK7wR7cWUn0pXlULiAIDFZqNEvaM7LmX4+5YQG9obF6
xZqu6LKzg2LMUI3fkc3XKY68TxQ3JPMCdZrKaunTLm8/kRYtCRL7k+nNVNeA9moq46fxz1oh+9ie
KCisAXBgjb5HqryDlRnZZ7h3HJEeaSlJKbsepmbyFsKy+XM6yAuKRLbJrFw3H9OvhYmRRA7pJcNZ
KBvK3CbjW5qQB9++2GYpe0p2Yu5pcDVjooC7OVk+4gnUvgppo34WmmGGahfePx5uxebNgX+e2+dl
rNbjlaZF/DQvf5kCxNEPZnNpV9mpA3odHZJS8BEQ0M6PQVhfeOsXZ2C6uwRG3Ca2qvAKIoYwEu+g
Oufe3tKvHCZ2eXLfVeHzRl84IqMd9UlM0YbBuWT4tP+LCfVvDqqHxETxP/NtrMQ+OlPy+iAHkdpf
nNDthw4+rOUtniDHs3BLnGFptnxnbvdTuAAr/TXWbtDsmeRnKBjmtWfIaUu/8IaRdJ3qEdXAXeGK
/93fI98SjZKJmqdnURm32nF1JmSmqnfpwsjhCv5/gMx5MDRQHS1W1t6t5iivux251bboh4bxOzks
G1u1JeGj5KKCmRyp6j8hScaFDIWJBgsvuCOw4rnxnBwPIJhi61BlUX7jwGXYLCevsGFKsTCqdAlS
Z5nE+S6fDTnbg7FTP7OcUb1xnjjqupv0fDOs0zMbRQtIM9Fa8t5/0gcBqvSjeqIu87ee5L9vqQN8
/iqoDIQDHMrK1pXa04Z7B7PSe8PTE5nEQkgQ7peBs0z2VFhax1tLUWBe/PJNKtEMbTFnLurdJZiL
dUzB0iCZQAfaDLA6U5xK2DJaSc1+5expoVuWbOPyFEkZXbmrX2ZZKiOq6VLkFYBbNAip8uHszmOV
bE9Aunam7b+6Vs2cCIU+TLsbybiz47u7SkjoqLfewHHCqCQknz/WLW4WN3LBNgQD88dkHS7HTfJl
SXOS+Q22mS3IaXRoOb2LQHe29Ufq2Vdb84Jp8WQEjRp32gQ3Hnu+0WCqgBufOrLHi2InkhwgQ656
rdovSKAlOrxve1pKUVNVwEMMDosOLPonM3jsVr9GHdrhGoWg5OvIuqkgx7HTPgo4WlS0QeXssbU4
JmtYrriWvV1ICFweoIgk0McOW+loVZU8i8KHOnkZEBsW7TwlCZgaQy1ilcmvbamP0t1gPiN+VMcf
EW5TITjsN8k8XRlukfSdsl0wGAgvHT5Th2FVqup3+fxLZ2ekin2UzlO518mDO2Ofyew8c4J6W4Y2
Wb3gQzoTQRoVhtKUDMaxvw1amKEIDD5Lo/FzyAvKD1HbG0e6KJDjXZXAG7s8mA2+zqPBzRxj+Lk4
Cdgwj5kwPLehUdDwGh030K1EMcbTFQbNNxR2JhuJHCWqKSYQG19tnOGM9J4p23rBeKoZtmaxOxMO
+p+GTdYdWmv9ACVWcmw9RF/UGbJLIvTrdY3ikT8pnmksnLdUjpg8IHoEfNaZwYJWPwY2Cv3BpkV2
K0POIgVw55OnAsRcAUd65Mq4CHenM0FiBnqSf7MlIvo3kLuReJ8RnD2P2kw+Ui2uxL2KYYy/1g4F
vw0efTneXXVq+4ttE0Y/fmS/se3tljL5+M+51WWzJZuo07mwCxiTxZ00cc9aueaoZzNatF5sq9z0
vcfuCD3P6FCTtriaKyHUcLuDM9ap0qBeHvKiCR+m5sZexK/0ivkvh7+rodL7K8P/gNB/gwI1IuTI
MDMfsg1p27ZCRPXCz/kvjq35guaFmINeBshbDagXIie2sJdGlP2cP2d8mOjJcnAgdydDvc8t0nZu
1LeRXX+Am/CQDAovS83SH+Cn+av07lwyTdAm9eQj3gpEvUoIaPbqdoQ2uXkHNybkHKbK09/bhIwC
kaJHQcfsGDQRYgTcTxX3a/G/OG5b1U4JHRP/N/hmhRCxHqSYEG3PMhJG6Zj6+7/floKaA1/SP0je
neibqMEbaMn6JIuRAQMuaE8BFyLNjgDJJmd0AkKoeapz0gxpqmZA/I9Kxl6D4tyrnM0V6c4lkMO9
7Dyi5r6Xln9RiN7JCro/7R3BuX5Yp2HqlLqi5JWYXN2Yjma90yvF0UwrPixVhUekeK8VhLKj1VFs
Dy1G4oSw7Kv1uG9+f5h0vFK/QRtoeOPKUsNqw3Ttyj3IuSvqHyvcEnhDUfJQJFr0/5N2O/Kl7ORX
9kSklPiAqtNwKra1LR/VkZYQXZwnFvbrBN0TVPpXvH+ASb2aBr4koJme6W2BEyR4swhMjzph5tNB
cRaCGqt7zNTlMEWUovl6TEOLznD6vpDl1hRcLhB/N0Se8wATK5BF/g8+2pLM2QEGob9TZW+4hQ7g
RvBHW66X78tkAgJLkf3sFlYsZ8TFX7SgiVQgHPamIShJM1gYVkCWPdChZxa2HKnz9WvULPw/CQNt
wQ7zXZ6lLjpV3KP8KSFI87vW6P1eJ9LRFSSDc1zrwBTCXm3K+1aOrgSyiHatbNFpcVcT9SlD700G
pWkruJyluGcOXsGP2IeDgya+Q5cu8B9SnGIfMChNB3mPrjJdxKCMyptfbI6q/fzBu7lYZWwX66Ui
+6xfzHtwz66VYUWlsvhBxz1D48tv/QZka4op+2M9il5d3rd2RWhn4+cUXpwznm8ThzrYnqyh2ukd
35ot2Dm9ZMWwiXd8z/MRolnvyf5tCCwnHbYdoorvid0I9B1LBgJD6iMoLgKwkRD1c0YCQF+OG7QY
ymZdtK/mq+0OEvOngGI5KuN8tNAOeHBOBovNB96BwbCz9MEyKa7m/PnXm+XZxEbx8LCDBd1AweL9
XnnNAaYTIKRL6yNxndeT/zc94QUFARhLLtoJgIhXyea21fhn8Ux+2on5gni13pMJ6ns9ObcDsxtK
STlbO2hFDv6e9/0mn48gNGNZ/MvtzjBtqAorIpQ9ZDbA247yUkPYbbXGwN0ElQFdrjvumqfU6Ovc
20wAYGI5A20vyFg0HAtBCLMnJlzioMku/aFkOdoxHSNZeIaqBhnMXGeISUIrWepGYA6ArBYk3iLU
EyrUXS8XYj6EJG7pZ0ejrbuGgrhVF5a4A08P8hLBNj9TYISCnjFlos1sEBVG4zrDQjFqBjT+aD0o
XrYSCDb8Sj81hRnpTI6qsSe2nG3JARsOwRr0dr8IhJOJcOOVfOvjkrb0Hf5K1xK8NatIZAdQuYVT
xtqDMxuIJfQHvSTEbRPXy57aZ/VE9gNu8UEiH0VRKnghi54SbmYSgZ9Zo0DVvKQLVK3UsfgYHu/U
dN7PDPoscFcT++U5KnpN+BTKVpmsAZwVriCIJHQtl2tbpcHcZ6Nxlp84Ern9EJ/DAOgV9h5a444D
5vk6s7jjY1QWVhGIcc10WKYMPw3mBfbakYZ47DXCYBpRrknq1m22cwBdhg0dsBoMsGHNaYKv2HVD
7xq7PpHTB5J+aEFiodQ3SkXyWo23OnkL3by1Xg7udH2IU64dN3jv0SaMANwpg8i3C0vyKYp+i9+o
3PJln253x5utLaIosdgtSENIT5G7HDJb3zvtNeZ8GnlWU693tGUIsuShyoWSj8wuaSUhER6kESeC
juTt0WdHD/yFWAw+gGUU4Zq7k2q+WuDhEOqD+9r7LDkkFaPjurEtLXVuB3GzXzEg72Hg9JiI8JGd
g0r2wdsdeem0cvey9jN9Zf+J9X9Yeke6lHVViT1QxONeT1cFdTLXd1JrmMll1Sl7ruLYCs9RJ49Z
RZrXpfBNMqfKiCxQ2pQiYTGgOAMbf/+Ge/y8laZw8Q5uxkUXQ/NEoyMjs8z9iPMiDb/G5siSNo7j
Juir3j5L+lzIx0RkpRuihHH75b5ZPPmCB/J62CID7LMU6eQ6OZqFhmaDichzxrozBWS5qq6HwcS+
Ato1zb3KJ7fxyiuF0l9mzgK/efXRMEiSpZrgCTj98KV7u18HN8RwI49GXvRQJR2J2KBc8o9Me2TX
OzKOPwc9LrmcxyJfwjPHpmFquLZLgyxPA36WpjhXuW8V+Mj5hpDiEmD+q8pJOkpKXa1QlHvMre06
iq3vrdj2s99Mw4OPpbTAVygDg74FdyRn7AjiXkYpihvoT0IdgpJFDLnp35x07ZtCB8A2XKHI7dLi
ApaLPbdy+JP8a1OIvzpkVdQRV51/GTwaEQnSPzvxkt60vjU28KWEwGq87+3Tt6qUOFiJdjHPE3Qu
ph70MUszhFHk+yjVQebSxr8wKBy8VNuSCtDqDiyCBPWszS9PACfqweycLcTlzyDbkYou8ug0kODi
DPlIgsRpXMrLSRp2c+1ZtTBg8KhEUECtT33CLBe3x/a64Tfjm9NZ9kbTQdwR2pi0pYqjLFsyzzPP
Qb60MIwL5qNKkYm3ZCvY1jenWWfxS9C1WT9/jR2weTupa8r3YbC+XUn94EuOwWAyAwmM6JCfA7Fs
dWz/v1gFel3dSt1rdZ/VgPz7tNCUpZbw2yEpn74PaSZAPr8d7U0vNPexu+F8DjMOwIeFECReKFiE
WXcL/M65sHZBCnBLMtYXUwLKrnW+WRRH9VGBA8PB4SsrZOJ0bNUJf+5AC2LFdyhiWRmD7rIPYaAG
B/YJs+RREsuvnfT31/kfPTAlNXxzSDRQtkqm9tqJLbiYVrlMgBfQeUxcqQZ02QbmoK2BKWcR4j47
omZFbO9EJbJQq+OHVZHT8i+SqVzb0TZTvU9JlNUbYy2wIN08Mpqducl0D10TXAIp0F9zEd7tESdO
OYbE4XxTv6AVUH9yW1hlDaB/+24ccqBl5Ia8vSIoO8AqMKuFHocjca5zubmQFfstn8GoVqAnGrs9
iBpZNfBR5qPDeCkC6ge/orvz+Btu5ddJj3LGJ34me+DwUKJq5WZuWxlEi5f2qebZ0LAg/Pvk/L7I
XnUgdU10wg3PzczhXJAycZnrTQs8XwdOW05TQbrNUVw1v8cqo8Rg82VMniJ7TNXHcvHQ2GkRVuj1
C5a94hVH/M6R8fIUdKEDUSr3erzRD3sG241mexgPUQ2/81gaBx0NHXuhNrRCG5Fxo9OXus1CdMoC
GFrnJSsgnS16EUbv0i7ZaVhDGEtWawI50Ow0ZsgyE4Bgz1nR+ijcQaSIrfxIUvNSbIfo6U2a0XIf
DttAwImvMs+371DM7XJHADrWzUmkp6QFUiFalKw4Z28pOLwoJs78Qq2qXzB0PtxK0zX0bNlZJMyA
PNO3S4UpDLTsgCX+ubuQhtxfFTq36mvIZKrBlZtJvmR1i9Pp9vdGXS2XWIqqiiqn+M3CPtkfQag3
56Ha846g7TiAlKOvfQ2HjnRFnAjstW/EFaJCqFGDLfUCv6exL1Bhiv35UhoFcNlwAZ/B1OjZd6AB
XXqNpwyxGXDX+hBzzCLyOKYJRW4sn6TzssC2VLFTSjc+FZwBhJu82MaM8cDh3hwfsA7Jc0oItKMb
prwuzqy4yILZRCez7QeOmwVZtOwtsdjm8n60JK5xMPvvFXeQT1gGun1tEYV3STZPU2SiYz5jJKBw
5FKP9aF97SWEg8jXpa+/nBXoS2tyH5FSC4Glbqns3HDJBI8I14w4zY1+Qg6TWp0KW20HJMb3O4F1
H8s0x7YfjZvkwMxwHzR9mKB5mt9XrdnEQoDSyVYivQC4oDz8OrJ2DAXhdwnteQZlZNA2UodeyiGM
ativTqLtohmev9N8JT1UukkPjbWdw2PuWxRj/NBBKjcgxrqWKh7qhismeb2LFQkUCOCYj3egxaK9
hlqzPxdnOcQvQMXs6TnksWm1sLo2SUd0McuVGpohLz2U+/ZmHIM/UCt9GRKLg2mL3+BOwhVtRIBI
abkCELFRy+6L2mXwYjnBSP0dV+I/LUdg8bkOXMuBDRL08mLutM/fRwjVX2PX/iQOa1Whk4yBWTHY
YLDK6geWSvvu7BrML/1aqoNPcCW85y45hcy9X7GJz5N2im32Vx1gWo6Kn2aU82vW3nbzxnzAYrp8
2X/gNFqvhRmK8cxZjjUx72D6xg6i96kLtm5nWuMyGSjHsMHtl6tKC66pAOXAy3iYLeW9WGkHoOSQ
833juoxRyi693kHiR/Ch0SzBNGjNnJX8u14Q6CwHsBiVudz6xrKT5yhK/dNHLKGfZS5Vn5zwz9Wz
N/QkbrksY6SG0HBbgbiwt0+TEh1Af46RODP6eqLxnMXj1q9H4DJ14dRbvq6oW2HKNccF6NDMTFXD
fSGjumFYfyDJQ7ajl1Ko9qiA8WzQ87NSZYPwt45znz1T7b+cxy+3Q/bgElvi9aUx2uKXo+BKjErj
FdquyPTp5q7mM+pdyl2fRtXn2CSoi6GUVaLEPKCuN9GqKSYRZNG6/gP3B3bEw1UJonuwH2EDq6+2
nHavAtZTCl5+clCzYTdzV/pvXXYKS3VaEsDIqsFTv3dMled1xSGJcAJ2g0n1L2tePBwp8sl7hgMy
rUCf4IwLyicpgYdZimsXIPG3RfwXBo5IIPbsCX6Qg7pVV273rq6M68AmqRT1rekW142zRwbr0Kd2
6p7iay7vOE0inlYNZbEcUXuSgTu40PpcgKcM3sisRfK01UYlfzOEaSrHfpQWkDdvFbViUyFfBKHM
0KWB04lQMXvI8pIVHS4xjV/VVg3j7z524YUIt76FlO/E2kqiCM8Dubieqdnx34s7NM4vT6D26UON
ieodDpRJWyxBSwQhVkHLmfcqD4gzmljFeFAEfOfPyz4dC7HuMpjU/ig53mp5fGeJBW2OjbL3gKRm
4ghILYd6t6WQBg33jCWDYWvY/7x6qoJmDjTGJJbxv3DJwvM+ok5m8lJQb9VrHVaAxFbx83wQx+ho
tznpSriXjrxEUessVIbTxgZP1I2xPApOAAW9nbbpT99kIu9wTBF+vlPhaoU0RnomJwWimWorutFg
+d6yZLaqeMomiZ0ypWvJBJxHCob2Whqs08mir2fskPCeQ1l/GHpRdt2bcpcT1N9EwGf28ORwylzE
9CWHyYdpT/hvbwOvKCyaERR75l/FdpdAPYmimyroqYh4+JFS1ul6NvVio6Yv8Vl9YNMjgYmPJQwB
gXOEv3FbHJvnGla3OecVH1Bay+JOP9MuxEa+4sPSdK2FE2dxTHvOdU/j3L0wHhJGsKxNzMpy/sde
Go1PhaDjvBwQgNPbHfI+1sUWX69Cce5dPeQmGLT9vkXtwaixJAIy7TuxypUNmVLN8gkxek9w291j
+7D2aBzeyxnYS9msdpOoyVeErdUDJCVNUY9FJEQCRWke7veHE2L2dS58cDf1uy07PCzbb51bsLyz
vu4fZK+aDL2fDEC17snJn8Dggk1EWkRiJpvn/N5hQSBllbCcmCvcP8FN17E31o5FUjC75zehKTFW
11OFToPPvHcl7j0XNvzEIg9ot98EIpJIMxj4KhPa5Ob+LogM+r4P895QdXLqk3I8SyHwGJx5Xuv2
ihglS4Vi1MmSTHhwcmrpPKPj9WODRC+2K6dkyj22tQIU4uHzUwvZXWjdcxyg8F3f8vlR02NA0Wlp
gswLq5vlv5xpxi5Okhq1EusAcS8SjbfGeYOUB0jvHsk8PTCNktz5qdsUfQo7AjGyo8YjcwQiFGVt
Yehmkf1szFy/3D33rtjDbXycEZgIw+XEORe5FVGDStuScBh+l7NW4s4ZN3MWVjusPF2EqhIXyael
r0yzDus73KnTwuDr3g8cOj/5A2uXdkjfYt7FBsuQI72OjyUsgChUs78uAfosfZHFVC5slFLZhgSU
QY8Z8BGuwg+m1MojVwwayU+npx1GTcLXXtl/VXz1cfVtz2VFiH7GSktMDV4QMhxtp+P6FuVrF1fk
ONwxhGun+wQiLitWyP+32IDy1lduxe0HOKaKTCUpNDNCyW5SxyAqhHHtuYnWQNqO8E8POEXA11OM
zUoS6PogZ+KJdsnyiwNvWrtLvRjfvYuIM2CDX4RH3QqjNziwiAT+YeQoc8UE0AMmnTyQ5ptPVJH+
tXfTVp8QdgVinA6HnZWKkjvah+zNyVhjrFUw+FY+dTiRtRhc64NNXseFIzhk/wC/UZk7I9xSyIQA
WxuaYEVBtPktJp+UYc2PrvgxG1754i1Jirt6A4DYZx0SPAmXZuCIIYM4QuqyDVall477cQb4S7LD
NsVAl+Lm5V48aOlBqsSmWYnUF+l0+8nBHh5nfwrPH8Wuw+ySbfyJ2zX2y8buTElnLgNIUQk3iEma
mTHqJEPxsRNJ0NCY/zAqIcqCo2PjlCj6KtQZxS5bWxH/crHxL9wyaAht0LLttDlkpTgXjoK8ZRfQ
DtnPU1uKRJWX/Na4AjarxbArQWYEeISWrzONto1dC+WeJA3jRdJ0XDE6h9VfKA3qVd+3RQ7M62d0
6hxTo3lyLZH/BPTnuRuA/HEjO4T5cNxhgrRei+ClmkrsRt25oWSqlyyAOk7Zl25aG6BA2S9s4Nn/
GqbQ7G1M8EmZ/gUAhSQF2v1yrf/2LBq7/zSM9IcG2Cy0DGx2ISC0Xngxeo40G6x6hTtdCDp2ZJWu
J8CBOQv9ZbqkVLPcCVKgykp7uRXCyhaJLSRDksnagPG/r6mNsdzqf1vbguBM69AgdMMRsEF9pMsT
aNQV5E05P9oWg4DsMLJjweQ7ZWyd6wA6WrxaXjSDrgwFJZgp+Y3PGFPddMcWiV5+msKonQLDDHYs
1lA0CGZ1pJoQon8TQCf7q3aV4THR4Ow2R3OW2BmxoG7wtZuxradONnftb3uyu4/50cMaascku39j
AyVl2h1/QVHB64vUtezjjc0JnKCtya3Aa3TCpUzChWz/A9cgRlzIucm3flMDVrUSAJ7WTEvYCWyt
MjmXZteH4Y/+qPYgzf/Vg9jlDp84QLMKXGpRqTSS1cu+T1VR/SjvF/6eQqWHRnJz1f6msdNPQags
Si2RRw2AF/bRCafvCtobdhWmnDEXoAcicejTT3DDKFO0O5oaBVT2KHX4q7G519kTUZuTjfCnaDAp
R9ZNuW1Qv+MaFO1H0n0IFEVYQ4KsYlnpl2ixk1IF7uVZiON0L8e2EHAg/rEF68fUTCArnhfqeI0z
rQoYX4PqG5843BP5L++NSTSKFey05ogoYHSC3nYVzquFc2zSfFL+gp7xVOVBpnyoQrZaBJkVrxoL
ofkbe/3gFd5NsRHcQ2I/ANpVYJgfRthCGHJ45YoLAcRNvM3PQMSH2cMX6zUArfEU3Q5iP00w8qaT
87iXv/h4kRnlH1zIdsXJDI7xYBDiUJmkzW9bB9cwVWhbj4MnUEnIPXpOPhCUBaT6YTL5z5JDywxh
QeNqFFho4zRoIiJoBf6YEMGmIyRr3ihGloG4ygsOEM8DqeQL262UmtKtsbsTY8gxjpU/wFz1jxZ9
WQsV91m1d3FSBdixPMtk3tzIbbigc6X4v6V1TKtQwrvI4s/IryxTnEWrGvnPprSBtDufIKzHwCNl
35wOcNFJEzwucjq0iOvxxOj6EhfVtjYvHLLjlmUdWQNyF86K6bcMXvBRrUpCqNBOsKmA1AfUb8g/
FZyVNaDTE78JOpq4b2bN7Hq70aPVO2cIBJ3uLPk2w5TRULl5q4Vqlo/By2/Pe+k/EuSvFSU0iLkJ
fp9988JbtivAqmb8Uwyl8/9YhEuT/gdRk8PMOfdiTe1j3ophdeLPNapMDkh7E1ka3/Sxv2K6gP0e
cQuJ9U0XeEhL1TtLSckxHLeln5u0osoL08A5DnjjYzwfxpA+kW1JLLaptxzxh+CTsm58ormp54D8
ScN95mjlvLQgpQ+c3kCP7VUS4hsFm5/JSxCTduapM4kki0otnEzSC9Lsbj+RHTdNjkiVI15gORyA
Hcy8LNej877j0hitasb6fPX67ePjH13dkrbTyDugwExZqTTzbOqVIPc2NJtpE/GRTkt1ZbFf0/CH
8TGKxC9BVPOQvXydm9F9EIZNb3RVLLnaSxpSTQVHhkYYLLD64J6c0bTMqGb29ECkMPD8iN+P0nIt
ufJqIvV1NzOlIG1DJ6NhZ8mtoEPUVraRwDN72gSojZrJJfPysPGCMyplQ/oyxBxTzSBaMECJGjmg
0zfwHaq3MYnRQfdmYsvAuYYuQBzSRY+mKY6kRz2b2bJyNrhIwCrys4j93UOzroR8NXT3PpoWgt2t
I/IEdLl+zLsoSmIMyjtvAJAl3zgMH/dgCXWlfaABDtRiZkGYBeHH4UTuSv8chRXKgixnHn98wUyr
4xBhNIA5DmMiOs6jl5GqXLrk2swlgDCBYk4D33K9CnBvki2OVQpH20wkDRsXicXtBYm2P4afUUIM
gQu+HmdtEkT53c3j2ERZD4JFmuwhlX5djAe3x9Grc/Q94Mv1gZOtKK7hL2CJoBizC+96SNc9vsR2
p9oQP7ECo//mi9repEKyxstVq0Ja7YRvfPicAQS2NqIsYQFwqkMHSQ+3aT4wBmLcovABQBANirhi
zcyvrfRXrnIpKEfcEi3JH1feONSa67qp5qbeyUBWpuvS9uLZAh2V7/Pg/zSB5NaVKQzu2x4DI7/3
c7JkP38cLdJq3kYYrvur9uQT8UVv73tiqg/iQ0WZsQBH3UsI9194gsnpluHL7eZfncPcKoC80s7a
Ioqsbs8EYK/7+q+nyB3O7beAatQBi97GWgGE8/O0i2ItL1gKo2t91VkJoWuP6pu5W9SJSla+lrKi
u0R/cOSnYAJZGFjBkmtiyjJsd/1/kwCBz4jxVE55esLW4fwHI5k/qnkgO8etjBa+SVzHmgigG6w3
nzLVDy/VKnwpeOhyUujmhfoQVqGqVoaW8ht8wnQ7UK5qj1MyQPAgpUVJwod+9hbJgNEHSlanbANk
7rDPFY6T8ZnQEHgukA6D9fiZNY3iDpdXWy103QckTntdC0oVqKc9N9UB7YkitFlWX/P1ChF2g+7d
/D1xzp9hPFz4WOkq05h9vxAZe0NSMuJjbFk38PFisy4bV4BKXsIsOSlwYWrxMyJs5334ofsYylS5
LJu3hdIHhLyLgVhJHa6R7V0NBRc4mzCeS/rNaYhmrG9vnO4bJzbbrnthE/d6Z9LPcL4m/dHG0dkH
wPOLLwUg3ikWp+lR5nza6HwFgs+ITqHnGY63OwhQ9M6FPHLi98pNpMezJW8MhYUILMv8kyxt+VLy
2/yuHIh8tSixKcgxZ7Dhw0tHdPMLRtpyAQ5POMqnT/+6DbP5TkqPDEhrlbA2ODZAQCpJrL5m7R/q
x8GUmf6DcoPBxHDZKJhgAid0C0mUmN3qqvwTKi8188GggQ8zsbewWhPiyNlw8YUfDKg9AK+q9b/N
LcX/hHQrXbGMns+oQS7Ej10ffL+C873bwvPsmQ2goVM9oTdDoCPtn7FmEXtXRCialC3vCsRDHmxm
LmVWveSUcEFYKUG74OLH0UPG5Bg7ye90Ww2PmolxIWOMEc9WPu+M1ERnFGm1lOgd/eq9MRFe6qWW
9qGnxXpB1MdPEhuV/P+rr8fo7JQKwHQvBv+ARAQiWmXvkViv79miNL+eBREsOCXb5noSkTuHuEsV
n/4fijoO0kxP+5FXl7WvJY7zLdMMN12Arqqy6rkCU1+mRHuQUlOFjr3N8c1/cTIfgiJBXPgqeylk
qx/lHNkzWTbUerDwBqGTHBl73Ruzb0zqdemuIE5OdP8jMJo53+aYFeuOOIxVJfG9moOxSa3KX1ru
MeRCmdBfTQqY/ZzSggoyHTRrzPdaDKDlHGnftWQcPAnzJNillicftWmdL8cT6auu8+UNk0BWzCtH
nL82GTrtOf6epxgrQc+kggT5j5zX0JSjYIUNzdpggh8UppQ2vLuVNaOvu2ZpA2J6V8wy6oBl2CCh
WqVB3Ds+fSPe/4fbDIEd27zmTRLZ3bqXX3dD5kRS2kow0JcFhh1E+VeN9AIROix2ST01zpm4ajs7
8bEs7lczdD2ZJHlux85pwuQrkZV6vBPmSOz1274eVSHJw6BLJCtO3AKiu0DiPGBg0a5tGMQhszLe
HC5K39bbTszwkNG8YAkuWhS3a/UQfma+Fbg9JFeOllFkez3B9VwTW8X+s2BrMEdnmTDdJ2Hiuwbz
uN/tZXtuykwfTpiNWEw23Pxpx1jI9cfn6xZdOlBymmU77lzYtgddz1R1R3XGU5Vgj1SDb4T6xkkj
CcMSlQA5vhkv9DE5brx9iuZbyh+53vqviiOp8JuzeJ9HccprK5TycAufWTGGQeYzhQ2XZ8FpcHUI
EguGWoJU452ndmx/uiuONSRkKVEvD3qVAuXJE2HThNuR64Azy0WibLeC0xsTwmBBdtqC7aTxHC1q
IoGiaAmlhpMVowqhFA9+k1nH0GNXKYmVjm9Y54LX3yiUllzbWZGJk7FIu+U/O/inzwYPe1CJMD+w
abDLgnunxuMIiX1z2wn8gpHJDOkYL1+ZKGAaBYoENfQD7pYNIwAv+GSllK/Zy1IZN1kJUIelMVEp
dxcpk0g0f0QQ1rT2UyDZOrofg+ShB9jacm+Hjs4Oh3bsy2s3VqiFvoEQ+UWcQa1bc55p2kwET+xg
FkedfvyKAOui89n9ResDmgAL9ElE4IU3nbPg5YH933JPUIwe5tPQOMbt4qq1P9+wHmT8vTMSkkDP
ABJPaR9kkOhi4RSsnkLC5/Za+O+wkAYDfepaQge//XEvJEWIP+yZm11JcEkgNWmwYLUmBjW/YncA
s8MA4xTIG5EjACGRLaOqnmqWRdaZ1Ye0cSi6cDwNKQFatNZjftbbKoPZTpB3SrdY7bLGak4nopGl
W8FZ6ImqX5EB/9rLPhX5UrmBkNXTtGD++FRjf5hYklieBeYDmknR3gXL9OAuJu/10555SNl7zb8j
J5m3faEvPSOe14CZdg8CmyhjGlbGnh6ugsYhdW2ejYapuW5WBjTlySogRVyyFS+SK6I0nTOUYMCK
rlv7heIJYAJfby8fYmAg6oju5l9J44+lg4+I3tz+kMEsZ73yKLt2+qM+ZPj5eAXyrYvwuNY3qPk9
rvGtt3hzav8OOcsQPOCgcO58ImAsRd0w5ojas75gIw4968CHVKBjNp6h8i/zzUIFhGkDPnZNmXYG
Wgpjl8Z3/GAZf22z6Xiify3abwbPvQKOawsoFopJ8pZMNEY5teuQeTxm0y7ygj1TQ1oMw+FOygwi
WtYckHYqN1z/oQg5Wig3ior02HTTUO9x6VLNjwEHc47HcCeOAXjM5XG8JsHBPYT+xpUgFh3on5mo
nHNsRPm4NBeUZrUjH0Dq2euUSZRJm7C4BBxEsgXEhoryalV0c91hMZWNDqlsQbw1LEfp6LIT+hcv
tTWkt7+ojjk4gu6llgIuKb2ghYUP52AFAbDrmmbdZLUkSdHdthIn3nVonEYC+iE5lx+eNDsMrtjS
HdJKv836c8Emj9zISHAAx6thUtJgFEJoOEZO8fXQ9JD7itjDY3PmvkJvpAFrI3Y5dfv2+gO0Vrku
Tfyyxvf3Y1e9eYwKUknA9FTQruifMaUtsU0znh/h7xELVgC18Il8zxVaCmAPFK0xtzYvqXQJNZIA
3oJVNIsPZ3t4BIPpEsxSaJGqGEhQIWOIuPxy+xksAX0x2P2KOMdmprvhFityTsLZQvknJjbNb55D
GRviA/ZDAacyqfdeIhl+JBSKyWDAJlc3uteAjXdYyY1czwo3lItRP9Be3ymjKVF2ZxLReT891kt9
Asu7clSubX+qv3UdadeVz8GE6GMkgFMh7THdiC3h3r9lrXwAThuB9hI8FmDOC1c0zWiVZnRQ3rHN
kS9LjI5BIShVXWQFL6kEuS1lZE+vrnTEqms+DncQ4R/Wh85HeYAOH+si+l3UgkGlCH2xb5Zzdk+o
8lvT/RA37b5ITcr0ENViFfqNFjRsSjGRiNjkaaft1tDXw6zxHUFrlnOKSsChRk8dor7VCLb+NGY6
JlIM5sDmkU62+izcud0AnPTG+azoWyzFAH0sueUKKvfLGkf7M1fPCIic3GoArOwaw4yxXvXPZYjl
sxaQEC9jaajk4wl8sHvTALaSi8CI1uxf57aymGQ5oe0+1q3DBsuCFdjHz2R6BPxXpe0bYHaetNDH
s7vEw7grMStshwQb+WVYCczCKBHyqQmuhJ8uYZ0GO3GbeXVtlXJ1/jd+Ae4Eum+wbxxw8ZRdYyD9
aGfTY8rZvy2Gi6S9LdJHOomQwylIV9C89kB2pfbse8gGOZdh6M1OHKb+fRClsyIS11mUi0zkYFvQ
vcrmpP8NXHTh8YKn2ARENtfnL+Sz7SwtzGNIqSxOCvGhbLeEDFH/wf9R2ez7Asji1ThKkZYT7o/O
alASi09eGNfAVgpYaChFmY/6u4dcU0kcn9EbmdzI9PzYM9V7tFuAVfRVS9CQ/MBHzuGiq3YE1iwp
aXmqRDllPQf+Or/6S/9j6aGlBq0CLMjcwUG0S6045bhRiz1D6Oo5fnr2OIALJ3mg70//jVCio+Dc
x42gRoq2bO/a+DW6YbGJoyA3OHGBHTPdnRLPuzC7pHe6A4ZKNSC+YIG7Ct7WIMmH5AC90e4Bhs6X
BsY5HF9k5//704J+m8+rnsRwWiQOQ8tbVjMXYV2cn7GQCCcSbg82q2zLbpRRBBSCabaCoeF9Qc+I
q54xOCewxxryaEncJVzmz1CSBr5lGjkIBMtdXjX04UrxO6CS4XG+Bb956CWt5Skt9cpkEwwVap7F
o/joAqRM3b8I4zZVf6Xl8T+3RLKcF/2OscQa0Ad0TzTxgK37uPOoUbyD8G92aX/FcTpSNIYO5nV4
c1o+76fzyGQc5Lcb0Tk3NWZxefJ5/sFOstURWlNi7Taoprw7zyvwx9rYFw+0ceg1rjGVtLt/tZj2
lQ5GstXmo7vMIB/295kWF13gx0M6GLLkK0fzAmT4fli59kB+E93HUrHzX1YbZDmmKiilGK5uDQD0
KHsnMvzR6Bdiyy7JP0PtZE8z5LV9oFBe7eli58oPG+W6zwGBbsiO1qsAUIr19QLvci0xSbhcgaP4
mAaFvcfwjkCkhKQZZXKXVYAvaKg93y4eXgXg920MKJZNcaWsJ34zFqSmV8zgxjzS2n4uYIOrvuo0
lsELLZgRoPVat/WhQq5Lu7WXCXg8uIIFhg7EVWJiCZU4Zlgkjl+bN3UXy1ELHIIXH1kFpGPLDkPx
bU68qsuYuMZKgBQOe27gb2OZg3c7ZvluE0BYIQESlYGF9hT62fSW08o52lcc+IILE3DkL25RB/ng
LByTnScfOfGPdagLLzRu2oK5mlANVph91Rqp3pD42o9/w2v53B5XdZz70/pq5mZS1iWI4C+Z7ORg
sdQwFwOTsawbJ0/jDEnyNlkO1YPbRyvuOoLlPdIgNxPr9aQAtAS8xlzFV/t/wncXiVw4WlaM4Cwy
wDf4pGFSp7tTEo5ajqSVV5RC5qFar9FhldwI6cF4fS7qWn93OpVmvpi7B5ytYs0PE5KvLvv4NiR0
i02k9jxbbOB0QOZ+E/tPIQOwd+JQwDdAAn7FFK7x5l2eM2I0Yz4TipBLNCiSjSdBlRawBEEUxohV
k9LFVI6rv9N+ovIWdm+6F5exSGekc86M6JQcxolFKJNmuJZhdXkK8/vrLQD+k8ZZl6Wg5lAM4C06
Psd0eLsn52a220hjnkWYJnjRIf6A3lx64IKg7H2Nm0g3u/NJ7d84NOixL3ZcDsosVo8z7/LsKwJh
Ie3gCmdzzlGM64hTyYHWnhmFE1an30ODybjJtCqocn0CjT994CUVgXB+tu2foK7R0P5Cw59BF0gr
6FpvXXh+A5WkxV2ZODvhZa67sh59srYgW1upjXbpjTxkrLX45QR3oy4Uf3DHW9vdfKJzdq230ip+
KCMB89pnOdGaH/mWSsL5ufq49eQedGQqIYi8/dKA2GeIQM4TcSoBEIoYLcYWza/2DXRfOhA1foEv
JLtUG9S1GL2BlicW5LqI23ILWLE9HOlV8TOHkr+ppECQFCIUtcgCDt9SS5r5DVScPohlauN2vEAJ
kWsKzT2o47F8r5e6KiTdefPJnlQ0vEjd48AzatMvKSvur/Z5/7GlzdavLGTHJJ/kDFaNSLpN6nFa
YQ/4+VOMn6WziwPpNqzQLKOl07jHUhUffU6OP+AQoIeDCx84MUF/qH4X03WqVp5/l/TdIJKzwkgA
rpa22mw3wdsY9DMWtu5QC1dGXIZ5wAHn5vzCutjsDpXE3eK7A8HRz3fNUzN78Vr63ytgt4ds8fF3
mCDqMyRro2KDGNTLz3Xr5PeYhmib8e/AbfmPXXEopOXxV6r6jrOtuvWOkMNjVVep/3Fq9V2e503i
Ug7oBFIM9h/10f8ipA0a+1ma/x2IcvLH9eFt1MNzCOkEOhtXehQ69L5Wd0FG0JmUz/EPR8JUjwYE
61yMSlYK/dw6TfPLlCKpEWrQqNXcWcikIaySyFDcMqNxYwY0w7lD0Ni92o8FK1p/Rw/+5Z2uvXjh
eZzZIby/lFYWEH5qNCo/F3egsFu1HuFc/7xYuGMlDpILe2VwogKXztzWI/iWGET7FGPUnb8GwxBd
qyHv8vpOk6jazPIJctX0dAnktF7rRk0ZFq+1IBWaN6k3SeOXAEF59GwPFfVyKTG6l06DupgKp3NC
F0n2iZ0czo3mOBu1hnrhCdMQSNIZ9cs3YW4m9MqKkfvT4forDJEdM09j74+71eCYvSrI11EExViw
40okaYBqUWp7onlva1BFs4c8u5rroQa0rq3eLMpN+SQr6oamOZgD4GudXe7hq7IswU4WW7HnqlAu
2jq20vb2p28R1yIn+v0fwzj653DfDEhlxt0ix0xF8V8Glycou/sOfvUCUFIKdB553Hflwv/LmHc4
ToUGVTgnfgKhGemEdHWcn+6gg2Qf4AJWfSxaCDEEAX/EwzX+Ez04TAE4cNI0A0MMJkefxwcIWUw+
GHblbQjcJocEAhhm2s+IRAoJnx5p51MHT7nFsIhJPyM2BNIKqxXIRTW/qChrGMAqBdFsgHTDag0L
ntdm6XHRoFIt57/2fAhW4k5iFVbO0VwafY2bWGmtlV6EKVstUX0LAq4XHp3jlRDQDkbemWuIv4sd
gvpEUQ+jS6TahUkt/czywgAj3mKJIUbixpKqU8OrvGzikGnrSihFurnHzPGaNZHlT8NTqhCx7FAQ
9iJaLFDw5tIktBQY/zmTM+lhKEZf2GnA7GFKgIXFjWxCP9bCzIecH03N6OGYX03EcTFjKUEW7mTv
pr70BFb+9s4kRqnDsR4g95u5dE50WVnnt1+4ehJ+v6mXEEyVpCk6qR8hrqBqwNBXMHk/FKzf0WYG
EfOUH8e/y9BZlPFDJljKPsGzH/PfrpyEi1qvZYyjzoASwFZ2omOdmJLpJyPw6NyBRoTaYXLqNtlA
CJdPDc2EHMIr1IVQ0Vxu6gQfBqJVFtPO6ccH6f/2Muo+RbQZ3AL+7Y18f/MpprSs4gUmgTp4TA3E
HraimTjQYLyTZe0k5wYODtHp8ZpsEI93YOtcr445NXQpyy+cJmEOhJE23wcNLkYIUEFOtZmXWbkf
cP22JQNzGdkYSNwr2I8H12r4eH1psXaVNgopZNUcnHPaf0ZiTNvMRM7xmDE8k2uJhSLiCxF3bayP
GMDXwZH33Hd3JxyvId/YCEp0CbR6nmewxa7dsn6ZvAgO/45cCV6b2sDj4EIRk4qFBtVWpLlDvk1Z
SBz+qzFti92SZmp1Sfg6ulHRvJtGOTm5Grvh6FYHKf8UJwRW6GYMNIZe6o0C7lqK7cRndy9L/EdK
htMsYeR41NdsNFhZzbUXDiumog+BQYmRf0PhoD/hDb9IodlfwRCIzyfj5tZadV2kBThXTuXbcvWf
fshIxNh+P1W/KRZVM28LUqqk4edBnBwC5gi9Y+FjsSQBIRDkmJkz3+ZnVakDpOALXjcu2sVT7hc8
RiVgiCtbY+eP3+TBuP2JqYMcVKQlTQSyoKYN6S+nvVkbD8VCFMJYA67BmK026LyS/X3OTDbFxq82
WjBZbLkDDkwY4K4Ok++hsIxq4nP90+wy9AvSWOkU8U4KmoOJpttG1In8O0xpDog/Wy3nUj0DzLgh
AHTb+bTILqhpUKmsIM3qzJ6Ps8uT+kkaNd4zmXpZIczDhQ77TaN2PFebcEK7s5XtESGM1WHUBXJ8
6EV/W4VwTwpeaSjhPmbG7uUUixufzwAaxawJCP0LwPkFrGN7ByMtfa8NfITDU7lEf352aHZX/uX7
6c2UVt3+DfSst8Z7CCUMcF1sfk9wvvvLobdRlqBamjyBuZZ5tjGt9nabPI7gBemT1fjDH5YkIKTY
CKb2qOtCVcH5OS7lJ4KWOJoagMcXx5sdNo85cH3h/N8hgbFmeEr1iWUbKlSbd2VUOmrElvQk30Mb
Kp52qYkHjgrRdeIIq9KAnyerEyJo2/lh4JYyPS04ikJG+6MXrXgi2mGiApNuY53sM8UjPOvXrsAT
O3y318A6E4pCXeHlwht+x7Fh3XKfIHtQS1DzVPHINxUqwbKwTo3Z7LJFWzTkMTZU3Al/MBLRl0Kg
30yoVSVh7neuJUwPWUh63olN8cwUL0s8ISBtyiVnj+wDW9yZfncimcvDQ+KixDGjQR0sH9nMyoLE
SEHN8rjpxypIDTyN38RQ3fy1IoAPJTC0XEIUDLQTffotF5ffy4qVXZtDBO66wycunnbzd7DuID5n
akhN7BjoSr6De9zYXmpS35AMfgDcddjhcSw6HES5py+SaWcZBNbvuV6OnR+dKmrShXqQcJi3niqX
Z/m8ZZVlZju9FdWZft7b3kS+wHxYhpN3ZdV/YxnXO2KA0m5E+qSv2JNi1SEKbgoNbSe+Upqqnum0
+5zZoEb9W4FOeqir3dAcvumulJEF7R83XMIOwh8JY/O4H4FO5UgyecZpkFQowTShAcJfsFRYe+Ad
My+ZHNgd9FgF3tyRe8ru+mZnkIeK/IY0/Bfg8UW8lxI5kaOfuQce1rKFvHtn5bk5Z36SORTwuR7F
bqa6C0dhJHFm0IBi6bI2zv+iVxAeFO5t05vB1f15teK/Hh9QyBVvskDlXBERzXqXo6QBadba/0mo
AmmP0+ELZHvjmOnagEo6Jqb39RHjgySE5mHq3acwJoudOQF022Ev5H6fJhn/2k6ORaY9BbdaZLIR
HSPdtNVzHJHTfTYZo/TF+KtMKdY85zK4TvGlk/eSCRcUvHsGe/hmqk3dsdlvMIsB4wgPmSnqipRI
P0lwqrlD3hFKJ/kSOuZ2o2UL5g5XGxMcP+ojwQd+uIk2o4M3cqX/8mYqHw3h+/Nyae7Ml46K/nzc
3H23Za9xUden+GON9tMNcj2MQlrtW9D4UVGx6fd+XOBcTml6im1N6B9t2/Uc5rsQbcNMsLxuUJcz
eqrhsHEMHX+GAh2P1XccOp/t6qz3EMiIn0bn9Tz5NRMumlRlqku5eoXlEHGZY1gVeuy7FhiZlSWx
sxWi1Obj87OfLgQETvqIEWDoexrUrJrvpk0NuH3nGiLuM3lXJSMzI6GEIN2tp3gD7uGtujetPmLI
Jq+N1k8ATcyotMrS6yKdIa3FOcyrLyotP/q0liXQuPciM/0+azuD0nIsWFCu3r7jQDl6nO9JwnBX
QmaZ0f4eAaVby9up/GIBmfbTORGSizW0j0un8IoDfPk2XH7C9EqsSqfCMimvO4kT18hiJG66LcvB
kPf0lSa3DPchZwxiiDSsFGLGaun0dcGxfd6ZuUNiwDrCDlXmV9q0+LiVl1G78SHNB02B59aiTIBa
aeKPRf9QMNknQD6tinkOH8F6IXttOG5t2ZXMhOaCaLU1yIZPLaLctJgy18XeMStNx6j+F/bd7mZE
XHCWZEYR8ao/KdrvXpaX3Tl+6yRpT/kgojfYQca6v2YNd5dyN+4FlftBuT7zInuTTqD10SvBkWNU
d1RDLspPH1yLV3TXoZ+Kyf5o/pgU83YG1YgDwwxp7koqW29XcLH0ZsPiQfFk0SvYrTv5nY6iS42Y
vDcYLPSsxmvpI67uKMdOCRnryCE3rZVtJUL/mAedQf6OGFArc5a43wjz8GmR64JZfwvOmVSnjQVt
E/bVi5BeFuUNoCBgSJkgAHSvg9B/SpNsPAGqzTGjDMuq8Tsn+swveCyRo+y1FGFdJrxNRX2QbsDr
1IpA2hckzH4gh72IdaFkZMksy8cIwZbFe/bpPSbzKFOvXWIhX0r4YIff9w4Ns0ggxcqQMnmrzLv1
OM8CEmZdz2nzjs9cux78S3Or27jnrG/1DOExylaobtZQr/MKTK7Pe0GHlRo1Pwy4ogtCKJBqYYAD
raDVPjEsogRErHXq8bSWH7rg9Lv13zuqHOrro/Hvfg43UvNEM4BjANzMlMDMHBxRWmQ+n+58T6ls
j27qveDjQcH3ips5aAShRgVGZIm3V9ea2I0t2mrYnhn2FD6Ky6E6yYgSJR/euMe+BB7odWhHxvQp
rgMGqwCQG3oGgbimunoGagqMPwhuELJcXQx24RIb01jNY1uGumWHJ/kM0ibxWnZy3nE4Mf7bobrX
J2mzLvokgAq4KSD6r4e7B1UxDSQ0+eFLoRYITERsYmVPNxmGPsmxb/u5vfWlgOWriuu5jBWDhYrD
UodGjbn25XOvKmubKLJh7OFnYFWaYfSqgZ1VjHqUcbYnhdmaleqzhSvnaD/jZYHLk6fBITn9SMLP
b5EmmcBGHRHT0zZU8fRnBk5p/v+6w3pmlSWy51RDhwqHCQAPnGaUCALx1GdViiX2531w5io0h7Ce
F/ht2w6dRMp724xk3Fhwxq+u09iLl30Ebze1YThjONz9YkgFX8S0TGjN5OJr+zjnYy6gOFt7gybw
Z6+3h+NtZLXgSSQprx7JVdUB4xXhyZ5osP4J/CWH4uTBvxR9lVfWw65WQYHcht52ZldR9zpfP5gS
PSKQ1jyjRMgt+RVa+u6jtBVowC7CxA40if3YEcX8E/+XIupWlBi8EZ+eObFwi/bEvA6p83VeAv7c
tNQXjCFfmCZ1RFO7SigWIfiuVvlFwT8QGRW/TMjdVcskX2xLJk0Hwzi8+B5FMYux96sMKOt+B7lQ
leRN46BzYLXIBE3buMw8UVWSbHNDGcn6gt0DRYMRIVu4E/y1pWDcwRh65AT8un0imBVwg02Fogbj
0IVBy9eQzke+2C/CNvR0hT02fBOw7Q+5uYb97Cg7LhAm7fxBwwM6LJznHYxLe7EyREQprD0PHx4f
t6Z1Kcv56puMxy9+BTlpjwUnYr0vBHnvvXrRSbUuzoPqO3D5yd81LP8UgB0C+HdOLCsfdtKYdZrY
1R2w2qWt0Zl2H7FLss5dvBjrihe8QQYISHaX3+8RGluwLMiCnDjwLbx8CQtepY974AC3BHPBKAvd
UYCnE65TmRGaEiQ0rdRfojlzWS3XdVISiBI5RoBxNfCBDW7foT7d8hR7heU6uOnLBu58vpErpD2G
9qt/XYaRHnn2LjepIkHuOGuoPtZwYQ02OR6To/G0IFguX99tORUJmRV5NAgMVfgN1YdNMEjz7JtQ
UZj6okGUBtJ/31guXFInV3BgpcmarCxiCjwtDOvRYNkDDNAUufoYfA6dpl+qhWyJEBTc6i6LsWip
kAJCu4MSwbW5XryGclJvt1mdS1El9YOjF11NqSvPxGtLXRTuGDSMuEvQtHx7avhQidGnYIJiGNtF
CZfxSl+YK9ZuZFQR99mr760OskKPoncK6dBi+pkzpSJeXQJBisL/pTZwkEv8pyNvwUkVEVg3svwq
OG9QQq9+awSoCymb3qwRlGJ5O5FU2tRxa2DYH8XOgGmw+9zFOPbHp0bCkH37S6VhiTaVG7SSDAYt
dKtpcDrclXeVr6jFWd7u4d8zqGUjJUcivjPBdg8t4Hgq7QBuWPdEjAvAivoClZrfVt8fD9uj/hJa
zY6IR3uxSg+gWxnt8esuZwqIXYtTBgCIPtknMcAjZ/8L1E7zOjk7ttSaHAqmBAJEkZMg7vSJIR7b
l4UOpjgn3wnv5itywnZRcgEhaSH0keWN66d3hB57JltBIoMvDbCPunkQblZdNwlPRfur/zTRyA2v
8q4oCCEXWGflch9FnFhcrkTmHRteCLQTqqH7TJzfvHcEJHl1TOKIe1Ddz9lVkDTh5HSWU9Lwji0B
49KKJw6FbdlCVrVH9wNQStHvJZwdUCYDg4lDMZsB+ABVI2gGl311dSXRf26cU+HV6K6V60V4Vkll
PqekxrMeGvpY+XJ2Um2WYyv8XXSxTvZS3BwyySWsyh+ZQTMC6x6L2yUydvwrO2GZYS56DyeCL+hP
i/jVl6hLYPx5lud0WbsYl1neFJnXRSVN7hvR++nuNRcFRLr3Ho3ShSwlzwVQBdeK6fOWIzX0z6iA
LUWMu/2d6wczPcr08Zmr+FpC28dJDf+zxVAKBQsbZ9IQBS6LsEUiIlmDxUiCubTvRNFZWLIWf1Ys
BLNMyUwYeBWHhGS/CpuPFwXrwZlMs9UKScaTdjjlLb77oK0m1mhpHJ2BRoOZAxB9MIf5Fbn2gJCR
bSXGihDxDIzgeOSjLgnYQq4xBHgFolikna8Ytpp1rv3A8QShsRr2uu/c4T3hmTQLuhENEmqKG0tW
LI5e4CHEr9UQ1cQZBSnHY5orAJqc9gqN1hBdM6HJ6bPqNHoCsyOihFdij9JQIE8MyiVkb3tf2SkI
unY37PgUFeks8pWxSU44ATP43dKoG0q++ZuNeMtMcRmyV3GUatH18hh3D81qOZ8ukhbRK+3N+Rbo
Oy5TfY8fQ//3cxG6bsXNxfcUL8DsYhXED9ZgS8PpAISFoMOzBbjIqRpPyherloFYsRSIwUBtHhyi
QBcVDLKl4YDKEr5XD9QylwvsvLhSg55/4URrtTkTffxe90JLQLXPyMRN5OLoD5jbT0ciMAh0UMCb
vgrSlLkRtP8GsSZlghOnOL3eb8wWrAewAUbvmwQAToCaCekX9ju36Lnti41OLocR2c/EHIhS4xbs
hb6bO8ohrJsxWXIAiqZWWQpNINrFGrwzTgYf4t13P8INavRmbUNZC+Gi8FdUepU0vZX1DmG+oUo/
VcG5SfbC2+P8mkkz06yPbswsFqOJkplFArBgx/zSWYBQm6zdNgxT+1wo31CUMF30seuac5ujQWx6
+cwt5ffuXaVV3Y+WHPMXJy1ydGiu74ARXNcD4niWzqZ2UcYHmbgj7TbjSswiqxrfQHhSjHSXtNSQ
uFBSJ48caEEe8CciY8kvoj5piXoJziyIW+JmOx9bqX6e/Bu2fR0bjhAzIRAPg1OA+Dm4UAM41BvB
u2Y+dBL6JzdlwBxCJkPdhnL8A4DB1QKaBc9RGIOjqAtbIXy3WS///XCQsJwP/6cNASmi1Xlb48DU
PUH0MFwDeTfiZM8MPZk0ZzR5OT1DqxJyIdyfKgYehkkw6upapEeIYpcBUBuNmphUw5DPFmgFsUoE
B6Us+07rrh2usfm4BLxyP+ahNpBrqJTXu3qKu2SSdUFUibW5bKXL6EL/zwsT+IGP03r+hZjMHrm4
2Q/vLRoYiH/R2t1eIdsf+i7IBfFf/kWOS5bm/sv0i50ki/hJ60Bsd32CckEv7EDmBjc+6NA9N1xw
XjcKoDNNyGrz3ORjiO0WM44D7Rco9ZuZkU+qDLUFbgaDe/t+G892ly82GewzSM2CBt8CUGVEiBo8
Vt6/uKyHzLUBn20rXGXCJLMvO1HSis9yFOWlDiMzJ6agblf8jMz5um1jY9hkXUS5PDMJ9y4QY1uK
psCz02TML6UDvxFudq6OYqXLv/KRRMXy28eF2h6fekh1wM0Kk4vWN+HFzdo3gLzYa+pRlHHuVZCZ
uyIY4B7ZI5V8PSL1sVTQvpsqcZc9Bp4jRbew7vQqOA4lHnYUNddba97yzH7Vkuxde7n36dEsfofX
znwOVpsB95jUc2v7SX3NX+eeXZqaRi2SY8jOuWsbTbbPnSbISq9IFjw9FM+N6cryWcI+15J7qMjR
0ekjW01kJhvB8Ldebk714G14IBSAe6s0egc90u7JGRoQHPPd0a0cLftSzqmNtVGpyi0++ebvb47x
2GXxH79XKJyuuWRhBBX6zS5LajbknyqUvsdSU0UsN9Sptug3uxGTc8WXkP3NegIPfZKdIlJpDMV/
89xlaqxvomEf2qVrJu2S9bSJsSGDpwf0pcw8+2o+gyxsM6umKLWq5U38dqq4SgUNJelJv8MmKg84
MGiT2d5p04J4P5/WDWf2m6scDBnb6f9zDat4dy2pWhkcQo4nzgUc0ew9Nwmq4LrbYeFuJSHsd139
FG7naHQ13LAbFfdf9OlnbYF7Zg+3JxxauqW8f2p69kZrKbe+UHzA8DnqKDoJ7qfxArcoNR9iXHgx
QeBNMSQeqJdAYYmeKifQjQrmoGPXOwPlEgOmC3ql/6Ck9pdpaZmeguANFnheQJiAekFOUtGrJqjD
DWs46YUxfAcyy5QCbAV1Hyodk3kl/J/ssa/cpmAQXwSPO8Odjuztr+Cp6/TnVXpn3JWxVHzfJqb/
L0qD1YAMx+kQKWgLfd98yDqxVxoF2HomWNjwZH/A/RgVY8kJnvVA2QecyHQFIqct17YBh5iVoiWa
Q2I797XrhWPTrAgAntKdOLFDjwN10t2g2tnQyoHsCZyTWaU4IcGzhHSBQ2/SmV02ZR+HMmmyPOZ2
gWJzSiP6DKXlZAO0NuH85UUOG5ciX+WnW/BM0ji2hRaDmSsqpYwovVABbGkOtf3qG+XaVTfnXbpP
FW8npydQItl4HAT7Skqckkk8ev/npVcOOW3d9AdfD+jMAaYqQCkUwwQJbvSYRlZQ4gBH6NIkH+eV
T8H+9Cq55fx8D6RjhbkU0KFO1JSkUQGYNZGaihgjF6d3MHtfhhU+bM6V0B5RrPGHbbmAZxzdwPd7
qSmZ/IRZ+aKPXORnhZsCKksI3efwjsFQgCLbhb7QmLpI9mx/0ZPFHW/yLR/Zwx/ZwEdlrrOUfPKo
qtrXMPl86zoTW/266Sg41M+q7Q8k6apv8bfSIVbG1uXjXtBfyIkpAlW9rmrSlUvbdDcjl3M5I+nt
ZaxQ8YSG3VLeFwL94FuSEhd3hZ1hEnXSYB2EP18P17qBkLQ2lOHaCb9ZUtPZIcUL1t4i5Q+ooqVx
aBDVqxvdmGtofVs2TssarA+DZFzHVwxbV49mHqSGS4/muGayNwxc8bJxECl27xHU4xSyFRAKq07o
Te/5kmy1oyRk3CFnh8jvuGzQTs7HRGaRycQ97dQg5Ix0o8kyGkxGBrUJTLn3Z/vhHDE8BaobcD+I
fVSL4PjRsbB+SWXvM2AM93XrfFfgdOH2bOWGsYl5PFiaoGvYbYQc1Vx6XLZtuK1NpqC1Oc+j0uM/
CMrYpK7GLfLTDxdaOlHoQzRUUM/tJ+jrB2YJjrVTEPLrQLbq9Mhc+gdeiIy6r37RjXbvAfdgxh/1
7Cs+3smtSPKdLLJ1EwB0ynzBncc2yvDJn+Vvv0hUgmerMWJM75Zgkm0ptErhuXMcKIZw63T3PXQD
eD9eAu1SUwswRlfobwakAdyuc/o7bJ3ShNxqfyODxyPXkNtW+CTksh3Hv1tbheTzxUUlu3oDOV1/
mUvYbU9MEExu5M/CMTM+UAH66xygSFrkV6cU2x/9FgNhOKcBQ+9xyDCG5hVd2eQk3QQZRjnlgBYu
OULQ1j6YWM32g1ukvQ4ksKrpwGL0eWgE7GPL2VZURsISpzh68mbblpJ5EWeejTIBFq1UTlV0cs1g
mi0cJNkS9wqE6CbElzBeI1Ob6VycAKn95FEaoxfM0D0jiOOuNzAM2fZPb+e3x4YoVVrUXcJvJlNQ
BqgZ44ZG0rHq5iYGJ8/2/6n7jOg1jKAPhViZBNAoFmlGRNwKoyF6RcCGwCh/cEtziXpTC4yGCPwb
2G0AHQUlK48UlnGvqKismRT9qmdol8NdrTGOt2ih2wvdHlDOEKK7fERm7rn5+fwfqp5jTx7x5u9e
aV3iiu7XnqP/hMATeP4oqd5+5V+pCZjB8SD7KndjKPK3jwGFTOcGRXU7KRSV5XOkhkWBF30BYk2N
Keb1dD74jhcBRZnobipLWz1oFyjI/GCVbJsvW0xJFNMLRC//Gxi2K+CULEOQ5FoUk1DlPdIRRFmX
U//MxKrobvJpp+NnbwR+dL0AsonF/sPzlsLuoIuZCcHsaqtSxrP5vA+WbdWq4N+tomrH8RCjnHO1
0w+2xlWyavbJljg+oUjrp4Aa2zGW+dc4S4Br/U5ncuSW3L9HqlB2SmscAQ16WiRaYC6DDzTIT6cF
yPEJoz3fCX5IpMMLeDXX//+bf3pOgYx+R2/CtqEmG47m74fcHUNPb8weIOce5mzPk+HRspYUg/Zq
8fiWCbRz3lUsuHB8/PUXm9IqDEs3hcxDFxaJhj/utnY65jw+YYtSezZROSXfW1CpHarD+gX6r2lP
IsqRj8ut63tO87r82f8VCg+k51VhfoBiLP+UlbWg/Nf9mUBS6k1eOvd3XgfEdzEoJN5e4lYPZbAQ
6vLtmrTtifDJdFMSrm4wVZYGFSnOhA7aQsGd1VWdhtJ0gJPaQKFRtugfVaboDcqQGFLzRp5F2coE
wAYUJQ3soLaWY7Fepvg7Uk781lkejdQIcKJ5r42Ux2S3aB6F+95bTIL/JEc2UePK6CwWZdxXj5nu
yKTtYje3XNX1MI0kw+VovzRqr5E/OdyHZ6lcZXdbs+fmAVrIMxWZy8tVL1LTEpWFkgvKcBSGpiQC
xJuTicJ39eraZSk6jELmrwM49w4ghr9KAjMU2eb24+O99roMCWyFdg5gDLJc/c/FNimCDICfE5kS
4h6ID2wMlD3EV5ov7A1tEBCjLFB/UN4xqH03fbjjfG3Cse3rp45S13GXzqvwDvX1V8z+fGfEgAP1
Ln98ZQutlx9ITBqggUf9+qahO9HIkbeKG/y9AE9+DDiWKkRlgjNFPKAgrpg3fTLl05WojjRPhd73
FkRZ3ekzwvNQMAhR297FVEk8jtF39RcaHl+6mo+wiWODJEA4BBY7QIl22tycT9ZACf2rUyyyE/vf
QvhGbqa7fEyLlBCXX68uBSP0lYsdLkC2CAiztPiOzA01P86VYliDBXSBqMAh6Pwdzd2Q8IgdfLNr
nL8sVo/Ear+o7jcI5bGUmRuw6koaW6vVhKlMc76iC8qWZ5WbbEItrmsBb1t/CDZJTdAjPxE7Hzw6
23fwvTk6R/KB0ZJPXMtN6SKcha1KOLJMoS7jlbZnvpIsKgjUsaZ8qnrfuwBcNmtSrauA7yYb5Aac
A+Va+Pth9Zo5T61eqUobNB8FvilfwaPKmhpJd6XPad0FrjDZa8gnGwBdK0zC8NnQgSP279FZHwfI
Bw8E7EJlXQYs+Xh/15asOUaBqNIeFwU2Cy4ev57+h6V/RUggKAha3OPQ0y0EyNo04Ludayep7es+
Qge2ADJF55Gwe+vKojAZm7l/xij6r3uQHbQSaOfcbHiH8cYRs9LCytfEGNo57t1RQbm853Huw2Fp
Pn7KXppuEZCFFsLSxQjT/G5cjBIlytjyDq3nJSTK99409Ni7yNDhFE/+dFOXP/dmRra/V5mcx97Z
II+tJMSaPsNNQ/gHZ5wf+S5VvxRWfGV/u4G/+GTMxWQph+YJ4lKwpGRXd4J/+Kjj47kBTyWAo1+8
EOtYO9kHNYENB8U8IaqLxNw1R8msSuYydG9Gwr9VMD7JpTh36ahQHqP/bB3skUUbq3tyfE88Yoy1
KE4jYyLA7bsAuwQJ43rlOLInCIImG6beQgcKpHRQTDi0mApFUotILTwDbLDfAw+Adl/WusqITtgn
dBDnEWBsjx1Fs6viDbgmrXGhuD9c9Qye1/vwSQvkUDqwf5ey3eSjpB5Xww6IBRfpunqJ7fT6/PkQ
RgaMQkVr8JrCFxu8KqdRWrn3f1JtKP4LxJNZae+XcWZezymhWRYtxV8LGCOp7ot0ZK/4XvOgHRqk
yJLUuhKzuJKF9hpmpWtNfoslhlTdpnCixIBOQW9FQjg9H19i8T4N5/4Qc1ylbZyjVBjZGhQZU3rg
HOb9ZX1/ZAtTXtbwzDCYnm1erc2PgVSLXaGYc5r+Rb53Ef4/MfBcOwoWvg3lcUnTkWcKWx4fr4pt
NP//o7rBX6AGTV0lzHTedB/kPF3mDzIAStABa7S2kV55pyx498yr5WDjo3PXPapM6cM7qck1jbtR
UM8aj5wyOcdJvPmwPEEWrxUBGNGkXn5LeIfhdDODgN+EeqSlUTl46DxACwTG1q7u69cQACxkuTqk
QsoUyVS+9mVFMc71mjRAnVMbMmniBrH218eROUa8IArvqO/gdVEaUSHJzUq8HF+qVzf4sx0iovxB
B3NQNbkTrfR/wfs/1d8nO5LmsdB1Bd/oDSt3qEyVAqj02dy9mukc+YzbOKm1Djyd6jpWcSrVKN4q
yER0X+LbxfGaPRqHLp8/ER3AewJ05KsiWExzMYL8OAvt5sIcrfr/pm7O2DyzhxeLzx2uXtHYEi0r
wFGlMnwe1Hwsx2/xYlD8ocVxKBmtDw6a5zki+vn3DBRGc+wEBjZc2dqhqgzgJOw8AhS27yTcBzEa
p0B5gWHGq1Zjy4HxTNgP1OLKq27h9ErydUHfSwSm3+lO2WCJnsxLCVNWy3ULo0PeQWbSSmZ+Kaom
cuMUnV74rZxB8FNv7ykfv0alMMRiDnq7nJve1LdmOeL939Mj9OBF/r9I4wva+bjmQD8GBQiVeGxv
RsTvLlBkzLwlZcW4KDOHrkyZ5GSmuP7ruTLOrcFxKOGSXim4m7XpFDugXJlunpYPW7kdZHSIrOKh
eo5nmIh4+6+4m91Lx/EpdBUWKSzCzlF/di+7FPhS7m3uG615jsvwCPM0/+/yWn/WVOYpPnnIgpqr
QAdx3PztZMJqm3f+HCstnRhp6jWZuw0tcumztfLr9/DzxS6UbS6wnjR3OSt25QGNCJcpWaJfwJNK
xm0GcQqAOPbwymVPr0sM1Jke+y6PEv5pMcWhCCtd1o4kPPogoSOvWhzNKjojzoJcb+PTrsMDnLo9
wzZRKCUQAb6c/4NMG1P0BbslzpwROsy5hDPoQWbQmbaqmEV8n1IOqybgJm7fbhaMrb4N5QE/UVDN
UoMrdwCAMCwc8PAw9Rpq/MhSBHNCAbRWh+rc5kSSSq8qsBsmc1S/FMZG4ABNNsEdGZZRslDhYN91
zG8Hjq4qa7ybrixdc9ueC+nSDpmCOkoOlrEfVnutVU6/mcZJFGINy8gx7b4Etgr0iwLm3IjMCTys
JFtj02jxQ7tk9iRx0pFdESN0YO79HI4t8FBNPNETX1TMTnZb35tPurNqo2Hgac02vBS1N342I9Rh
Ts9V2FVqTA/vyHDBUIooWaCpl41RwriIH/hClmQPUH8QtHB0WCxlmcWPAnGr6f4bKEun+m/tdQyD
PukBu2ssT8VWtKE+1Tw294g22S6yRel6hREnEawtlcgE6aBkSCtoZuHRaQ4mhcKU220dHavEzlE0
hC/y0b8uoUrBik7OqkT7l+Dyy2xJQK/8xwj1I2xAZ2Xb+HWv3ePID7tjQCNVeD0luVL4HD7I9g6y
2DZqIrzYKOG49ynTpl364sw4Uo8AR6N9dp5ZkRgYZy1h9TgE9PFV7RIwdO1ixRXbotGP3Q982Z9J
t3eGGU2YPAFN8vmcduMXd49zLZYrDYMS23TnvmGZk3G4jUel/55e0df7MOyNGr393bK2izTCDCSe
f7bTGAal0c4GpY8+veN7tfVhU6IqyEwVyc1yOzYCxdQa1yznFQ2a5UEF+R+KPQitj4UPWB+yyIG4
q+12bGi/edPbgpXhzLDnGR6uUVUzRmWS/ZC4eM5EPAGgb4RF1/aO4dvlxy5r4Zss9tVa/0Qbv/gV
e4RneForwuoixny3HMpocNI7GOqTpHfdgurs/RJwP2YHwy4CHYJZ2yPwfmNsPXdKIaAvgPRK4/xx
LmiFvBm/+peN4XgUWh8kvGK2PY5sOin0SO0MBP3j/1Lti4F5JRtqoyzdjbOu+ztNGwkV/l1GHeMr
IW3CbYoTkNz2KGGzsj9gdEJgjfHyY22C8yJatkC4S59EhOkX9MjbT/9DRo0aLBB0xR3lT/57DO1e
iR7jjm5sgjnu2BPfBrZV+vmwYvhn76KMDX0/IZdHFQGpKwgYGTEnLFOmEv1EJqjmw26aqQ0DDg8y
04qoWZzyTbkBJbHu6kevw5BFnfP01OWAK7xkTliZL+IrxqFWhcYA+6/GuYsir2g8kpNtsglkhXfO
kYWfZNFc/UQCBXgBlULKCABzBNlK1NLHbYmaEFMvPD296LaLq39kmwKCfn+L4vd+ALDb7qOshEHE
+plXIz0CGhZA/IZRuCqqLF4vf1VGs+VeH0nmDPVYBkHp5/sfT0Mq2CjtPKwZ6fF04vWb+Is+p7/4
v088/NrvmygLDwp+WroeLQAZHnPigD8PkxurMXDKuM8HSyu/FBLKZwZloKPH9OqbT4YptgKj/DM2
H55U1fVNYpK7JF/wh00cWM6IbrKH+ynpJqpAfN86Tc54c2TdiMmZJQ0WwBWPD7xEAqbc1+Wa1HCS
60z09VEuxjJSTIq4eaWePEYvXRG4jKA0q/l7ON29rC8Q3+uiY2FDD58yinhyqjrrwrBLOIrOiBt3
qPjdvtvgBfISrEE/fn01aFHef6jIO3vsYCPm8XOsMij8tLFMbc3eLYtdsNXq9KrAfwOtXpZ0QD6J
SBwhew1pU+HuDRQxp1WlGBe6pSNW6WywYLAlyfJo2C0zajRW/DsyvsfYqk8NmetHfaUmTeezAhB1
v6rnZ1l7Df36eA/1uiSQKuRKpVW9yaYzJYTvFpR0xSDqZIxhnPWnDNsilWk3A8KCneXnGvxqHHuE
di+NBqUqbfUgV/SQFvD/0T021YXGeMg1K5U1j18hXLp82oPrR5vcbyyqsikw2p8M13neqPLeoq7R
IDtQqagvIPfxp7fRsPtkk+momNLfNk6KEbAAXGa5ej/yRuGiW2CLeJhlCmCwRcQRxFqAvhgXNFTh
IxQx5XLDvG4PIJ4hxLjEXZIqMJRfu/A5xe30GLTiE55dskAlAeM5DZxygOiLyOvEQ300JsQ2NAlf
zTO/YVby+IRA8Ao2JqR2eaAq5iQtvh6qFgm++ETDO8eTIf/uSqsxXsuRLfja2c8977YDbgyxlW9C
QBPCxPrX96ruqxyCiycSafsZha//TL7gBl73Ht5OKICJAp/d3v0Vd3+8rcRHCW9xDB/lYLaftcZ+
GmEPZVki8ELsJYdPFbRdBgI/QF657ijvGXIgFLG5wxNYRHA0vGNtdJQjQUZ/vix3nQDeclhij/QH
Jm6Zd0Dy1jYtWAEjqvVIX8zBb5ZFkmCyX4EVh5VWR8ngSess94ZGyb2UsLkX0WTOG5gxYfT0TFia
9OJsSe3ZfiaafEcfhY0vx6xmOmwbrx2SCYPHwRdxDTDZotqPhxKvgX6PYksS4nBlVllVjeeovMRs
xj46RNb39ecyH7dMbIKtcMCcARMNrfWkzqiFzpzbocLJp1rwUDwG5WEnrZNZpIe/G8SxrFaJV9a1
9L8PqcrBA6892Q/WFJFJa8Ell6DOGWdjN4oDVNsg/BDKIOINd5LfJEVpxL0/QpqpPFsmLMzQh9S7
GCXQyHGzcahHUqypMhzE7vac3AF/8fTcFPPWjMmG5nVkM+BgdkTC+2M78zbK3ucoLUBGOLeALJ9b
nA2czpaDXzrtcH3VLDEGgbJj13LJFuEP1u7U1t6Qi0+1mHXL43RrBka3t53sBmoe58uxlppIa2Jh
Dy2b6O9RunhR63i/53EZQ4f4DthkUclEai+BTcn98Auxubkmj1DJHa5vTjhps+7e1un9v6Z87+bf
NufnzXws4HM6T8ysm3gtIu/6MLXyVqxwZG+pEcjXJtH7pmtfJQiIKOhIjjJXa0zmKDyhXBBgC1zR
D3HAhRKAxL76jywdKrUXf66v5rWMsFcYoODBoiG8DJ+a78Af8I1A1sMtp0ccRTqWwBpiEuhULW2H
dkgI40s5G0UlrNz3u1Gw6qtTgVaUyi5bxUuBbvRjc5c+TKXhgCOKlrwa1XUoJg6EmibRcy6yDFz/
FC8rcJU/Ucb1G1uUYaUjIsMrhmWg4wdCI+1CJAyEu0hI4Y3om/nFGCcvdxC7quViiDDeO/zTIw8P
tqRMOdfy424JrSb4lb6TbwlphWIuje5s+42bW7hqIIIBOP8mLYgAmLl7nFdN/PCmBRzEC0NsH3TI
W9Yvo+U6PYqdfPZPnWKgYLi/vGPqNoILCUF73QrtZ9wgO+vnR/4yPYolKz5324hO0bKMM728Vp0+
Nv5poqMpCezgmyrKHQQkD9W3e3RE3GZBrXSF59gjejDH7bNCXlPFJtx5LQPTsosBCWKU9R+KyTIH
fXWis+UHXLGocEYqAkF4mWNoO0XH4j3S7N+f34PdtnUsDX22NXd7/hVQA9hk0dt3P6XnbPcn53xv
PqZQ+ghE/aYiTE9wFaz1ckDlxXoEWsWq+x/XJh2oUQuWP9V5X4Fi54AeWaos/qH+BUk13w/2bR7O
tNK9T/2GvvuJVrM0G2CpjC2vFSKuMad/fWsSzHoNJ9Mg66N05NHjjxQBs0w0E9sECEcsF+g7mrtt
mJ+6F0Ii6AIRLsBKvawL7IlJ/RxbU6AWMJMDnT8bMvI3FP3RGI+74z343e7yzlLMMQHvwFNsCjP5
sPH4wdJ1EKtaElgBateBUApt5AJBJBNMk3hzMfF/T0zl9bK6CxyCe8oYvho5GxxUNKgSG4ZkE2K+
eHjxDUBWXGTZMvwwEWzrp1Ghz+64yDFJ/Y97+0MV3eBd2HgPIAYDUJk4Ra2MdEmecLAl+2g0XDDt
X/AgEQxrPcKcEi8Os6xu9iaS1eS/OaWb7rPKBaIhqd0skffKKZBpvgp0oBIJcmuZbydMg9G5erng
RTwrNQ7mpDA3NVUgwOXWUid9hcEF+xkohBRSZ9wyjk8ZFMkXNO0fPOXJQoqWUXFznhoW1Ok89Q7O
VtjTb7SeGfEipk8S93seKlXL17XrrLgW7SV9UHfaa0KhwcnbRt4Une/FYAPpyoB0eOxy2aKTD5SE
khF+fSqBifYDE/lUSoV3TEH5+J5jeL0iy5woKtkzU6BgnTnSxIcuLrgTRlRZYdkJHr7ZOCanCtWM
Q+fjpkwOqAFbLRhbSuRRXayNH+k10qjcs90vPkPUeOhRsxepT00rLPRUjdGXD7pnLtSslO4Z+mYu
ZLZgYis6VuSt/NtDYDgV6bN9RIs7F337NwZudR2O2WJ0EX+7J0cGziaZNXilcXrf+Do0JFLqZtUE
qT6Ku3mVf73S5QA5awLHykGX9XQaB3ie/qBGHY+alMndPuF8ypKafg8ZoCgmfwgJ5iPopbHArMjo
kt43t8WTGKIH+hph7ud1cR6KQ4dcIydTQx8n2MmAh11S9Taw8jZH44yGtgT2Hl6kMxts0R19Nyvn
l52ilUmiHZ3y3k2FkZf/KFERImpcvLNEF/t3gwLnBxS95LpFXHPezq3CvPtS7RclmPSPBmrQm+e+
5Y+qjCAO43NFLpMMDMIGZtfz0VKmU0gDl8QpI1i22I+Jb1c94UhzWIwaZK0UjC2gXHKMQw+eHTq/
iYfsXGKtZ3N0Pu91vK1GuMuJ/NJ9kvM9mLlVC8rId1oR7JR7dPRqxoCmfnvoo2m1uH8pj/HIzsE4
HaUApVzXmKZRMfQiN1oA/lL8dKwUsUMa3xP1PMW6Lr/hyQZTqf3wz23p+QnlSxSGvvCx8RTWh/3U
2RvRX+A2IyQuOGZJZuutwKG8W+FKAkDvXoT45R3yr9jbqXfqxnz+nICL9MRt+4mBThiIkCWjhzV5
3EA4o+fy6ihgzFB32Z9jb7r3QUqaMZlMowCxOPBTdQbFZGDxNVBUJLAWp6XSUnklAwb18iiyC10n
I5BDKiIk4/gv1hdNKx3fQt8iVLIu37JnGAiZXox1FaOhtha7a5JpDRzffoDk2zhOIzxPqBaLO7U2
eIskAitF5bBljLX9NnG+I0mFnrQzCmSwqZK7Q8/Z/nDVMwzqFKuBiBqitqF9v5hFrq7eC5l6a21D
NvOfUm8nGiucZLH3zsAh/UKywNwbw/cxBHlOGpVQbREJLV8GMhGWqTpIShBIqwX+OfLahgCmJRU0
96lxKoEWIiKC04Re7YHTHKkbWxhwYEw+rSYgOnhxPM8SBEOsw5NiJVbe9I6FIJjkcdnVzpxfb5v8
S0tWy0qpOWRz5VusOy9z/TPIYvUfANjFvN80WyFXuUchij7mX6ixJ4Cx6IvjNBXoZchw2PG12Tro
kUIO4e0ZlgluoqYjFpTTIRw/CwzLnlTbtZCrO5vj1kSKcYyv2XKv+kR/pbpuSIFoicHKaKuotMva
WSoW5A5TXNuhKHRV9p6knn2eTmQIRUjP/2uhpFrV2oNTzckZx70N1p1iut2dnEHb9yEN3IploSMD
laEiaIgqO09yLfOUkr5iUD2mgJdawGadOlVbJuyC9cdp+YKgryBepy/S1+XBBf1r/lUJcBiVmAAq
mdTzncdgmx+4nMz2SKyd+xFDXvwqW39AJAI5dc5yAdEqFFSGv/lCKnNobfn/ROuOX5Ek4f7uB7TC
xDYwZdfKzaDCJ2ypbhrL6EBtRTMhQcUp2ik3cNlHRUoQWntPM+ZyTOY6C7JdQcwsWlEdNrD6tJPH
aHQSS2fl/piLA8Xr0XolcO/B9DedIlSqBzgS0tJwKhbxAjrJbgQiuIaHLActPuJRO6qB8BwLFP3V
NSrVnvJdLdCZ5CEGLvyVFcaIm8yO1AX9UtTfjAGderPm74YdP5Km4CWt2DbWsqKp4+RC4yXec5AW
zv/0cdZTBLjl16nIm7UXoDK10gcXCu6V4ZbHv8/gDG4VqvBWiFhi1ppPrN25XSwsY5zFsv0r6NFT
09h7WrfjOW+yC9PFT9EDaZu8j9L2AnBcFdgbFC8o7saSbyvb3L+xzNnFS3XqbeBwqp1OmX4S7WmS
Md3m+XN3TXNMp98h+h5jFJc184Wmf1LY7as6sU70/kB79TDxk+ZkYMhl00HIy8EZvZtjzAcZEk/8
3F/cBnCVlxOcey3taB8QeZFmLX89pmcfxI5rsoCP8iCYKv5GcUUb5o2rqLXMRI9fsJ9eA4hITlNp
u0OLdncVim9RhRZK8yJaDpD9ZuOQGPoc9DBe8qCYcZp9+hFQQGjlYs9u21Nquhi9l3DgzuKXyDfz
rmos7qjNddRsP2Brhr8b2HeyddKzW032gIqz6JRQKqQ+n3GkZAAnOMcHq3/n+HHG11m2FmpSUE6f
Ss+Vuvy45c8RDkTQEQ1LczQKrV2vXRfTnu4AvxqsSM0ET3RyCHuUTUbXdSrNh7zZ8czNhc6URLbP
yEE4+dJkspSfY7hu/A6Pb+vXz/q0Wcc9VbRstVOrsL3jbjULGpVIqpAHDJ3CVtk+vKQUONF0O6T8
lwBcsI+6gmM9t2FOotY+oZFPlREOPOEoh2Z8JsHl5biZpMcasq5g3XjNfJZNIHhuIPENi+du7mA+
kGZ6xg1B0E01GFiv4qp4HOo7frBjHRphio3SvQioNv9tx2sCdZdkGp/NdzRDBIy4egE4R5DGwO1c
EHGMvIwvG5Hepx+UnvsDlcRvkXmfOUFNr5/pb9WYo8p7U+oZ8cvgEOcWeM+RT6NB2iZzpNgfuMpx
noWC2o9TTysu+G17sqfuoWIfNlZ1b0IJbGNqu0QDCfswQHoGJq+ojI9Nnsr8t8OfHAaT5tgl6lz9
sVaDZxuT2LLrOF8hqUz/VNNn4KZItsLmLb4/AeMVZqj/NsUKYbxCmaHWFPezQv/mL4Hsdpuofksg
fDnmxkwISfftGN78p5aX1H/a+69/+muLQD8JoYuh+J7zFoMjJlVVDQHqS6lU/b+3fvVjAjGB5za7
n436JzV6pdN26SZeGcdi1Xqg21rRBvvdvmil5W3Jk1lRubyCaMWzVWG5IG+zYzXWkpRCg6eRorxk
o7neIXJy9f9cVbxIjxc7IH8wCul9N/+incAZliE8r24XhcY/1Ou90IY5m1aXh37XF/DeBG3wNnmm
VrsJZ3qP8naZTy7eSTt/J2rdxvfJHWhZ7haNOXYU3JZ6I6NasKk+pZA/+ea4owvcuh9NXbrCsSCf
TFLc7DQfsyd0Ac8AnBfohpL2iZHtgfut8z74upAF2CbkbrhIOmRMnPhfDeUVfyGa75hpbBi98FWP
qf2FFlGGtcINQqWWoiqSFayTe5spDyXaqS8HaY16bLTsQ7XLuwRlgiE7oqmkG/eABceTKK+9qfTb
8GCDV0VJlh6JhFKbmQoGcj+T9S5dOZkr6PN57x3zdFTJ9TFIwzgUIM2vPrEVXS46Ud+0hq9OLfCt
K1nI03w6O7elAOX7qAXN1IHEZW0FJEwvuyZjjFjP8iRjptcGOVjVyJfXIvOfPySi20ATOCUblDqi
ifXF8jmQnLOIfT1zzMLp8Fp9ocBrW78h8lA/eAnuIGdaySElkwlvdxVd2VFs3QkPVCqnGjpEYYAq
J2Bp73kHIuvA5as/psxfmRAbefThGw2B7Gm55xWkei7k6JK1NuZAD0kJ9htYaS+wA8xzY8ReTO2X
vi+PzPwh1l5CxfssFiCsmowkvtSDjvOTR7R4NowG8MKw/sDL/Oo8sswYpK766DP9A4f3ti1ND+w0
cuM05LtKTE71VwCf1rQNpL7uKhLg1AUh7cK6NEEB8kOzNB44FmE/HebJVPqGfkNfcMJvRw+ozSNy
dIaX5jbp/jVy3eLHrTrMwSh2EuSd6sF9i2EvRYkaD8qdOcm7w57MLF4rKNJqyigc+1r6D/BpF5tS
cXM3BGxRfj3LTl/W8g9nq6tf2cBPvbtyYckbxWmA7NnnTdlgn2illMjt7L7NxUjVaDaxqMe7gUNF
9aFl750Cjxevm73YRcYUCLfvAd0FNsZ54vn/WjG5ugJfic6qwUe9hQMGROFMBJHtB8BnNkGfdHaU
pIWJX5YgzuxgfDpxLJt4lEtN6f1/wtEP2pHcQP4OPmEqhPjA01ztCrvmRNsOGVjgokDYnKd+V4QI
ISPr+++pKSE3P6zcLlSLV6x5Yj9XREs71Xa+JhMwUXEDV7M2BW261PLYDgST1yQgbMDa5rcvshYW
feNRrmrSwKRzGVNhs9Q4Wj99YqNqqDc33NKNw/yJsZ/rldQLWzkj3bbQoiLEDvdEnFBEllCRHh4F
AAaiWPT59fcK9HFgBuExBrzX3BZe4ecDV2tSj4/H+TrJYVdiA9y/WpXAtxUpyc17pRsGDraNXl7W
L/AicccVddJwmwDtm78P3BSIofnSBy6WsLH4isFnjq1DEEMyZjVzcorCTdVaCmh21SnjmK2LkOYJ
OQHge8NJqokb846EbGfUco95M9T8ieklxrxQWfAABb8kAAeLlpTr0eBukxdO+x6EddEDOMbY8jDG
1lbusA+45tVndRViryHt1O+Q4ZAhOWBlpMyN/5vsHvGqQD/U7rBhV1pQRMFliIoZk0ADi7Ul82TY
tSyw1DTAT4eYxnTgzkbTvas5iYhZEcEbdHcZvkv5TPkkraSkjdP29X8XgQDnRPI987x/zKvZFbVU
LAOJkibXv9ZEY3G7mEMVnmyZi1t9qztAeNVd1LB7sz+WYg5NEA9+SuF9yBvMaXBqDExpAwTPfMlx
yDXgSngCWAXj1mDbSQ1DQFPaPxLI+rbz8SbNfjHBwbH/S7AIN91ZBxgdvUeMqQko+CCyC1UD3O5E
SPfIRiXWwySGanXuB5Qg/Nr8a+DMYaOKLwNgyda2hEDmvo0RFKRQXZcSmIDz85s0+5uTXRBr/O1I
OJ/An4psYjqANvx50+ZZ0PJRTWwRHJf00nwiD+3kZ5IWEzNNGqSHgnYlyoRT7/wMdU/dRbw8cIB5
TRjHvyxx2qbH62B/EjHySUP4kSfjNP/l246r4gd9WLfKH2BOHs6ieu3cqZXB0oQVDKmR4jVjeeE6
Stzty5/rNPu37mZbG1xF0K/QlHdI440SM88rLAWoguMDFl1Mq9FRjxUCzYS+K04k0iNJ3TRnKG/E
AvQQriqg1c3eUANIEKCFQ/e1OJ21XocA8U4A49iJeBHu8M+VytYul+Pqprem67oPpHKkbaxPkbxW
3boi3f6igb7Z1ezerttq7W3pSEnRgpnTZ5gBg67NynbG5JM/Dkt3iHqq4HRyNo4wE8eOllpxq0mC
OAQooebYZtqJZdvnT3Pa7+uG3u5wWRd93EJ8BrS6gsCqfjGmEfL4cELdldeY78YaWlk6/3OwSwYH
hM+D1jGCSQovIbWpvFYQZmJ9uGsKgrNprS52hXMiP8Q5u42XYKKK0tO5LVxuGBEcWrD+zNcyqHJm
C10JItV51HyIR+idxCXW91rdLpDijE49voZC7l3NFiq/ailVqCFTWN27nNJ3njr/Efy/7hxS2+EH
oGomirdg0+bcmYdk7P90mlW2qUrTrlzTQw5fDbcTJ7C8uFRuy5mqtY4/PFdHPqGBkkD0TR0TZ0K7
XDkcP9oR4mglma0/m2qGZKLGbVmDtmUNbE9bWloGfDRi/OBovcTHgPUXInFIWc+Gl+wAD/5X5w5G
v8KDgufnNaW6jNGPNyMwrZDtqBCSiLHw90cAfuq4OlFkT1AUaNknZCqDkidFb90QKR5rg4APKkLV
fYBQnJ9x+K1Ojui9kKZQ+9RTGsXPcDNdN28pF+Y63r916w1SWCg/dE3O7mirTDAgH+8cNv+3Lswd
2/65LSDtX6t77CQngs+Tl1YJvIFAKL3EZHML2yxC4Hgd/12PHk/KUx0/imJaRowqXJ+y5aFxTDq2
ypkxG2BVnF1/wJKkQ5u/GCVM/aim8UCw09QIOPZhcbQ88CZx8gXju5fb4z/Y2JIXVNEBfWl2vaGh
PygyGFptRtHd1n+wFEOISAtsNO2D1QPp6iNI0vBkGFr95mc1lZAjYpgItXnf/MRlaM7CQ+Vc2slw
X8h1a920tBd16IPTHFVA+TLXIr1E7MC/DjYKIZZUtgT7B6nk7wCiXv2Fsa7ndWWCmBYTXkpQG6ao
Yj/ljPXLhjscjGjkl4+U+ux//aUY5NWANb8XH1rVRt9hUits5or4TdbE6ciyTCQQ+lS/tMJRa9x8
F7oIvej7qt6PiJFu6kugTENhRacd+zflmQtey8/T1UG9iP8IOGK6u4t6BetVmKuzi/aau0Y+TbeS
ZCUp56jp/1Ak4/Pw8P0GWvGfWqMBosGv/tHcdUBKG6zYEWGf7PaINXO0A5UTosqlWQ98OoHld67I
PZ0DUP4Ds+jxisvZbmfTtj9EFmo4twcsUcN1qtBF7v/ScmRTZ/xgKARrw8B1DFSbjpXZ/6/Cxa5h
L0IZQqbdk1RDTsquIuNBhbmO75XSQ6Yj4NH0xUBvpR3lLu8bzxdumFvUZ9I/gONOOOBGKWfBiYbH
XqSVzeZCePNsPi7gfY58VWcIRqXo2+ZcyfZTf7Hp6waGduhG2906s3auAYFhXtCqVKyUrRV21c9o
32h6b5b1yEBUp1VzRVvanQwzlqxPfxEEjayGu1AzC8i2sWVkaHb/n//SWrgkCmF3n1RVc86rHu+V
9b2Jb5FJydsE96vYjRcTBR06jnXZc98hk07t69RaUfatyBEAeI5/TfSyRiev675YvZXPRnm2AsZN
JKO+Q/KVlJA+bdEhTzLE+U5nLxsk2adHVWkrcM0bO5p202ujGPg9o44L4dyu5YDfVTjSGMdFea/G
ZOGubUs1T5mWzatn63YrpRBPnWh6XKjwbuUv4pYx1/MmshjbUzlh+3X4qRey+xwN3fDTeETwN/Ml
LCUUKoTgiKwWWkNDIqzh1T186nZTsY46nnyEDNTsui0N6idGeQEm+GH3IV/dvfoEeSf8/gMaKIOR
lXd+/Mi3VtlHaw4dgoECPF/zwBtmzHtJ3xBZstVKw4Ncsg8LTPaBAk04zSTm3Ald4TeA3fVNBqDK
99WsOM/qflbi1A2QrDKS+tBuQHtFjOviDVOaU0kGUYcLlDwIc/npMTnP9oWp5hIu01Hjh9g/GN+s
yBc9b5cGGzaWSDcOXXqw8PycP0fu6GTHRzeCoB29PXrtlSUNZdP9+WQocMQ5CrSB6llrtAQ/UBRQ
HOIOm5fCG+ohue1yRupClDE905uPbztZ0o2a1kAxKqG88nHXQvwe/sIfxpk6AazH3pjHNT4//lOK
RCAHpERw53jjAapQtYZS3HMhXq7ovNxodCkv88skxWUwpPp2UWYp3YKrHs7OfZWHkCSlhL10bBDF
BVj8PrObo81jHjvKTyXIGb0l7NGdpFbZVuiBTCwyXaZEUf1V6KfqJWKnMyqdmgMVd5hLq7KlTojo
j3ChfdwmLiDrhAgwbL1M+PAaQTAgAfCvGhnIKFVRDY2IqCBxG9GU6Ot6ANA72LLdGmNn3IuQVmHu
uWFluD8QHhYHCePLQ7t7zEIa44rLpD0PrUqrQD0/vvgHUq35giaSiR11DsLhC+f3peinxbehF8Rb
G+dwciP+y8jq0yzxDwM/uTeIYPl+z1YETMy519y0k6Vy7M4OkE3DRwnfFggwSZdNy0bv2mIM1xka
9odnRIurAOuXsbOxp2/Ricg9/kofcza9/KjwwQXIssekh4LwvLXfv4P5lQHEQPhxOVMeE7SPQrIz
KzeRCRmu4AnfKR0Rn/NNrXYkgZnpO+tXX4MTNDpox1dNbs53eiuSYkgvuUO+z9KWNiL9yImAHIan
YhGr56IbD5eyV8XUruxcnpj6cacJflPwNDX2eddmvMNY/1BnDAN8z0QzixBn0w8rOSxyVRk2Ery0
tDj+AxADtFX01htsqjohQFv0vATDFJEr7tiwnKRXqmD6RSX/0ncllbe4gIVNErPi1EptZCspO1ny
9emXx787ruEdUxXRyIDCBFMnK9AzCUewlC79n1I6hj1d8XQTa1pobkus2Wm5nyrxcHl0lido1qPb
an43+Y2QJTIiE0igUki2Zjto1HCge2Icr7tYy18NelgD0/ifxK10xnpnOg5BVcw9Pe8irsD6c+hW
yL5jMZGZH0WOE8pR0sgt3bh0ieRbi8ffb1l+nqkURVZYwQ7VacINxamZfXgzHpLMN1+Q1EXaufrA
sMptc4egUCWSnISPxUdaQUoFwGkEtCH9GpPAwLUiGVKgopvGcXJBFvGmkM1dfwa2ANaJGdWQPD1F
a/zVcjAtAgGjTZWfroBW0p+Fom6xXg9hsRLhSkkl0/hYZc2bn1bumj9LPAr1AE56yhqdIykNWHdj
O8CM7FyB9bp+csvxk7B2uiJ4wY5ds0DRNYI9hF16xJoBHDJ+tIJXOPXloL5cNjKPwqgtQFwAFtWY
qbfhdzrjYFdJHF0SAhcKcnf4b4NAX0unFimk3DePw5qB7wKrfS+OZ/UIsUnjcWi/+p6fsQTtG8kS
JEq+B8o4lnXOYvY5yT/zI8dBgo0Hxgqem7SNih66GCFSA+YZHLECnCIgJNLBNjZQOLeVg2CNu9RQ
/D2aqeAyF09MmNT+BuGdqd8F9VfL+mjPMEeuwCc/ZUomSBETVIHW+1vzt6/dOZrLwS4llNcYegM9
CGr07MZv+6G/qrOnvYJDNqf9oPgwknzVvUlWokaE0KcEx5ql4fNezmlsoUVo7BLk5fZDIHTRoZb8
H41muGTpwo5A9p6PykVejKXzPr2ufWnJ8mPG+Uu2tu2ih0vOx2xCjxMPwGZStnQ3Weqjf8L3RvcS
EdymFvMAXFL7HX2dCcoTp4Tyt57h0z9+mBvBHllrMZ2ewsAlSjHb1KIbtXkVW4/in7nTy/4AlaKr
Sc+V+JlhP/ZNHCihOXeg3BA6+rb8oJDukegtRyvMs8UdvUbwY41CT08Txgw9a3ukRKrzIyu8E8Z3
fXZazjycwYGOTeQNMct7WXNiNRFqa1HDl6wlck2PKkUfNaGyYBeHnvNXnfbLlF22CFvCW0Xd8wMV
D0CgEoxnGuy8mGjo4BQz3B5nKMJ7yHeUXStO7u2iCEyd5+KTYLI6ZDMwT3GL4n+0C1LIPuWf7VgY
k84/iORxfhLzBAFQY6eX044XNFS/5z0+J5a51+Fv74Vpum9EdkrKWB5L0BM90kRtMZ/6xr6c3bc4
83oYJX2SuPaz04DnQaAfNuEQFs3flT2UnJ+zbBf78pX7/9yMKCoGt5GgN330L0OntJP9JKiLVfVc
2UdI507Jljl2DprKQ6XdAAri4jrZPCPL9iTMhQXUUJ4VoMU3bPyuZ9UKu3XAz8RIn7gnJPkw3GW4
VqV+ZVIq8zxtyQgD5NONg21vDHCmNJ1WMQcYUAdSQwBTV8d98wzYkTdCPyLFr7aX76POjX+ZxWWi
v80hw9583tjXGx6vPCvegzpUGFgflUsMhxb8UuagLeFNUw7+BXpKTGup4ktI6IRRC+gG6u8Fcama
MlXDzAxh6i53rVfoBWU3cmPGAv0nkL/aMPPXwxuQ37jvNn0X4RaHvQP2K0fZ6o1tgEg1jmou+ccb
MCCmRXG49zp6CB6R9aL/0EsMNEf5Kq48CsPXopNn97PrGVG+RZBk5GNjgoKsxcxbLXUDVxLjvuVu
Dcb556ijr62egVLmkD1n0RtbN137hG9VKydCvTsykNMLMdvEYxuY5uc+ed3a1aGP+RyGUWUUWnCl
DyFf1LlDmbqOOpS7lHyt1UA1eArg9xQJs10yxyNNLVsV/nLE0esrF6RERQNgiVGkjRIZUxspf/dd
q9cYcp1p3bafr4J9NOo984CGDCQfl3s8QEVKA52FY6Jr/QTnsVlRf/G1x2kLx4TYDwIeFodS55n6
aKC/ybk+jvDXkZUsRhbhpUoH8MYxX793pBcS6bkl/KoODGtZzyEcl2kdGzJFRTTYJUX4k4jr4sgo
i/sPM9pntE1Iomi1oaQDRFnSjwhyrfN1KbT9Es+ocRf9P+JnfwaEkgdGRVGd2KmIyHN9rujoXSwp
vfwdXfdeIuRtpqrw2xsx7Kij490CEWRg2oJaCXUmC0QqWrvub9etvKD0OsErOM48W/9h+UcCRKvd
8BzxsYRcsq6kiCxXm3+iPC3mqQ1xbZk/A8r/sfQ8nl9KLevyfWTNymX/KHPZrOKpyeGtpbo1llox
p2PPY0Ng5mWSEzda9mmKjafHU2q03ed64hClugM1HrvISxcU/HSAA/qN9r9yXaNbNxte1xYVplYo
BSpicQ6m+UzcxkYXI9PxNGcEk7Wg1PwuEk4uXy2WjoZTrtEI4TOixLywA6EyMBtkxR+zFJGHuL7S
m9XtaJVy1tlwmgP71gtd6WPd3l67xjOnCWlUT4S9oNYZZv9/hQnFbeep5NwbY/aIfdE2MlcrDg1w
21tidYm2dlM+nDcKThOGMNmBVSXmrPlvzfTr4bBd7eLaMp/KPJh0SWPxKkfzlN9mUfsUf5xJtP3w
em9pjQvJKgcZzR32PI7hKk/ysXiVW/xPAZklbarAC2YXhXvD5IUYPXnpq91yS/FgJxCW0sM8nyQm
R/ZDmJip19Ghx1lMtHxpJuVuKbeCVufZYbZowkOTyljysNhIuMEz4DwLFZI1WbottIqkQD9ETrET
L9plI/pTf112UEEXgAMUrk16q2gCUMrd3EVSsRkfNaPPsIYn76GscrcL7duoTL5Pf/zJH25Ym4xP
E2qiXLeyxlpIQeMfYMS9aerEtWLnP4zDHOUN9+f66I6BuysoxB7qqLiSM95YHb6hj4HdoGV+qxaq
ccEw/75yiaNBpd06m2z1trDbw255CMvbc4Jf+mqvNzLDJ3gVK4eCSJ/gQWSVi3PbdSwmeZUrAw4k
sSKo2sROY6c/ctKKk5kh8DXLm2E/fPl/lKiUr0kS4Tf2ShQY9LWypOcQ5Opkx3nKf0UobikX8PVq
CQQ484nngcXuolrRylYwFeb0G4QJwylQylzbED6lFuUTMgBFwgfbLCOoEije143DPdgY23b3r4UI
jcZPyDwWGGm3D0AZ9dQYa/ISr8kYN51U2EaQd0vY7hrU2k1zvvgr2JRGRUIicrXA8E4siNWQk2v4
RfEE7/o+hdO0yEJ9PTIQVT9NRqoY38hAv2n5KGos4aeV+c1Gfa87vfmW8Xml3wpPK/ddOv5YOoiT
jlsw/j+Ff0zSjZWCaImJE/KBsupttD6qWIKP44Ru8EcYo+XGhw/e9hlNEdTQ5ZEo18zQMwMXhbP0
TSAq2vSF2/XazTUpgZE/tu19SqXYuFpmKNiJyJY8DYsMfZSTL8135OGf7K3tIRJU1nDLI4TofNbZ
NTxKc40T4hmjLMqnuxqNVYno3hkSWPmqjt7qIzf7dDJGi6lfkfk6Uk4dIYUYtkZsKwKe5fLUt63W
QyUnUoUNVzWDQcKziqYaeo8irGEzi5AnlBfNEfKNWA+ejr0N120IHks90Mxo+AgMmmxrPs/uhjsz
0HW2NWwjpQbkSNQKERclq2iAGc1/4SZUAeITVd4Wa5PrzzRxzH6Ah4OWP1cWSICK7sUBcNy48lkp
NIRphhySqCFRZbsnhAUy5/ZkW2hdGCKt8xi08+cCngbYulo1WMEQAD+6ytrsT7+1xGqWhpI03qaw
X6KFVZnoTnVj0QIuxHEy600Jd0hmaWEmvo0jScCBlLNTqrkTwlljvVa5lpD8/uTW939AC2FVslyk
TEigSI44PiI90RBxoQ8ZGWcjU8dnmcEa3PjZJTGfJe0caLuFn/9s/WB5vg3Y8jgRrNC60GungOLX
h4fnSRJg55aX2ZU+UTWqc88chWY+z6fEIwthgDav/px85h9VtiL5c3QJM8uwDnIRIKGzfAgbBTpN
Xs02XBXjw8L9PklncIBXss2pN5Qu4oLrUSI4rRGNuBRhqcwp9860mBrviLncWRbGObZbHqlrILmd
6vf1QvhhlzSWRRhZzt3sNw6R+px83V408DBKtVx+LqQGggdpkOwl+lqYNKaACZpuKhznOLHpbTxn
ECBPjjttZcbjPgS4jB8CKYfzeSlWgF+xlVuDAgB4rt+XzGTfujZon98w0+H4iIZ4aMmfH/RRFtms
l8GUSNfSUJL4hHdKVsDUnwf7Ekz+OjntJab4QrB5zOB8doUzMODgyO8ItSs16lGbpaviuJWiEFwZ
JNv6Dv5iQuKaSJBm+QfN0CejLuCBiJehZzlGgDofwIe0L/FyVdAWOZnWnSYW7FZzNcU7xlLWTFgS
nTpgmzXCLoChnaZVnr3yGM7fsln/TSeDDMk1HGwXdU2oo2bzIja9huS7jnz2jMhT5oVcLXBOfxkB
8fa9J9YOZsuBWXLWAKlWJkZ6NlKwx6pIoyDRFBUYEcZvBULW4z/bYyBSOGebwVUtzpq1H96Dfg2A
hee4yW2h6C97F9L/UaHqYQwkOFhc7VOiFfvKugi5z4FXNrDcIY12oMKcP7LoB60+qv/+Ih9n+3lo
C4HXsL+AI/soAtOTmEzmKF9vOXP9kx5FcG9LekmdolLtBso31iCwL4Oyv1Xf5wffedQ2cpff/4tW
XMV6cjfqPAnlcfNWy2tNkD0tXZZUf2tUBD8ndJPo+ToqSeyaCcQ7aav1QDB66st1UTKYdHdcQw38
jyvHfS9TCmXMG2oABAp9bEirmrHfCBftRqub/tk5Cjp7pcsxbnBsSE5wJW7hXKgf59UqLbT51AGu
osHTT44BqxJoT3ndHnQPwdDelG+YS6QC4goHluF5yqKSiUD6vwu1dJZFKzYvqtB8QbDNPhJYB3lR
BmHnAMR+wEEqi+wYsFT6uy9jGYt944qPS5tWowIXEJwFleK819BEamQbMakJrztPRs8nrJ+2rO6+
HR+ekzdiSTACu72UTxu7bH3M4jPDemHSvHQ+ZJFSY+zEQadOrbw5NSazcoK9RHVU9RScgTRrxPk3
I1dPinZh5gA4DlNRA0Kk+JJq6wA+ukpphzIwdZVQg4VmqCE7AHxOu7foqDQtl8jOQm5hwajO9zJT
XJBwXmUcxwvCEdAjyvh3sefOercKvp6Tu2W6sAb3NlfqmGU6sOVZU8g2ardEWFakcA1j1tXeptDF
I5g4//pSJEHlUTH45wLNa4p1FUSUV3Nso5/uCgN7upfVkwMCrAz796jrwEIU+qwZpvU3aIbuiMql
ZgqRgxmXzkPM8f0OCxqsIuaGSRKUatsulw0pYSMyOmolUnTrS0ulTSO7PFDb9uJnvfWwTs8sIUoe
v6OIwHZVl6iH/pdQPfWEH7uncVJ+jgdLUEuA6rzscbRXuc57qZJGSlSSpM5YKZ7RUo52jZuUbHp3
kRbfSli7NYthVyFj2zgHZTkCDIBu8wG1mTry2M5SiMucdHcB/6x4JqbgpiU+SFGii+p2CBoLPpwd
2j7FPVVzQTQoOUcCX+lspEKIpRdtkWZ87bFQ4SttYI0zqwKkJVpO2p9OZnXiGaEIYUKfx746vXTS
xAYzg2pE+6mldLERM9tayiT6ymk4ffdeXRPYNRLt1ZQXvvLv0tZ+Sd23CybzSc5BZTjUSgwB8gjb
uWlQ5e2pZa9Kwmj1T/EmRO1wF8zhrLveM9LibruAVSluhaxiLO3b8uVnHpHlZZ9YECx4GNyO8OJf
nGfm6uvd2328MDVTKN5da4eAtkHNREd0KU9LMuMtbSrBuOwPtl0mEaoRwMsiBvXtiXHT2YRfjvy5
ZnbWLalcIrow1j3V7wBOVgmh+cymFk6o1TydLqlPlegUx0dzwr4N4WrtaNrLNwY8z+P/VSjSZiKs
V51aGJJa48vBvbx+5EuMl0vEhu2fiHUW3oMkQHlCfHddSXCH6JX8UAwuwkYl2uxbh4WzlZ30Zzms
2cW893K/UzlWa3sb71F97L6mqDLhI57a8FV1aVMSuMw46RZH0AkaCm1Ltpi4co+0KIY+W2UvDmSE
Wajt3UGZQReU8xzXTj3seBQ/ha+rnKMzi9zLwX86k3m0RdGYvMn3VU4rMPdk17eGteBx2FbuCp22
76nyEoYKhxvvk684dAvqEbEmQMhFIs9gnj3vLj8KEjD0qFZ7pNaeruGLiwJk9zKBkBaDz7DuUIZi
24rEVB4Vbi5mr9n0HLnF+THW6FxsixQXom6o4dkAf0I1+PMZnXwBG4vacl+zGkNO/b6/fiyLpdY1
HdRzUojTJTzbqtUk+P3NssYtgXs96ZYSZiAQCu1RswV0e9rpVmgKev7kx/NDZri6KnXXGGUDlrNT
saNK6eacTkqJ3034of3J7znsSZep6qB/euk+aM9L229bJKSZ7vESqHfNpoUu6gGHZ4fkiyD9bA8M
1GkfPDjS4BNbxMOeU2VRtSEtd+fayokc/uGNHiw1usXlf+ApPCDX9RljU/W3BRR8bQqCtKR/Y4XW
x5Rf7sHpwi3kWNPqa12kgNy6lWKXCRPGHbjbbLBco9BEIg5dKDn1Ss9xN6DEsOrVEqMoDP/Hl5cN
cMfgm1ASy8VxG7xQgQm9m7vM0Ewnt4rw9XUpf6/0Yx+cPxteLqgACcqylEO+22u6y9De24gpP0yF
AX+9MK1c4pV+HRzp+pO1nkcxDaUXpy2ljO6ge0WyucnwFaxdHVKZFVIj+WUg8c97/V/0I0uE5f54
yS7IzlZT/fEXIRwA89ogvFcUmpGNZMzw26ItdNMOSRf3Y9ATGRNq9Nic1Y28xoJqZsHUOnq1CY56
vneNIrpzXQrHCsTWjuzXF1LgsLb8umArcKSqAdXWgA5D1KOqcIQaKpX0TIPP9iH/zEJxnglOnxl+
N5mcVOtBo0RCnY8fChR5iwelz6emAKb5iYtp1AOinaeShqwubajgCnLNZdtdnq6jZXX3jE6MiIEB
80Eu4jOXPS3H7hnrd21FGlUs/3OW1NCwqOXuuxdegMYJcX3GooIa/prvZ5Ig9cz3Lykyp1DefV11
FtU/GUXDucAHUPwo9Cy2mKBnkK42hbVDoDEzYo1pX1U831WPFwJGn7KNWANbOJsU4l/63jQxJXA6
ozUKgcxsAgpLBo4say6W+0VhtMb9w8OWmyUfF8e5SsHv3kebsa+vHU0pA7DU5JjcuzBSvU0ldawr
3prQa++uhW7T3Enm2VrLHr8J+eFWGcWSltggTuhUekreNu2r4dcirQ8t5zQrnMBCe0ZWaV9DbZmG
SA8N/QVCxon9w6mPwYUFAOWYaKZbjiTG2Pv8wmkkHQeRO75F1YY/s2EFb7tWoGZ57ZiRxhDy/BgU
dVibvyPGrhutjZgSMyvfAz6kZv8HAM5XkkAovxzTHINM8iRDy4e063Fh0B0duO97krrP+tZCqj9E
Omw7nYMjIGJzFSE/Ts5m34H2IewomnyDU9bibGoDfn2hleD83dc9AZT7MArlg6vUx38oBYTQx8zj
jEYX/aZI/f1JNQjqgkYuWOIr4zTlIjBooQdjxnDGMhPY61y8kZOheYmLZ0xHSnziY0BphRfF/mse
cZv3Ul4jQNpUpVYsxZr243iWZopzkOTVRgQaSWLxoIrowVPMal1iU5jZtaaGe9SxPf2YDgqvG5NQ
ESm6dYFzu5g8KuQ5cIWg4+cAx+zMczx2VIeQDXIN0+0Tl7cc2SK9I+FYMqr9iadKMLBg4nYt4Mhk
3JqBjPWazb5UPt9Ksmk3ILqUCk0/g1VJoSs7HEcmQmRAh9uGWXzYOCtsOTFjBWSvNGr88NVwyG4n
hYmrLyshMGDpFrmw08Iz6BObxM6Dqqrq+puGnyhjgyhirfmWqDunwshfC9GwwrejQPyYiHUePCuD
Yz/ijrTNcxFDFFEEBSuu1wStPvN1i1GRERVIW8lkwRd1Wjn/0lA6cJ5+CwcwKOCrHE9ZMAHOSAzK
CA6VNSoqsHa8cGgELKC0NWpzVxFJwdKTfYRHy1RukMWLgamGGUHDt2A6ieaaq+YV/YQDUdNVI8Gi
feH45REtREudOClyT3C4K7S49WaNXs2wciflHOW8a8sMmLjHr4aF6hP3TOmVmtfRFxPr4+LmXv10
ULyVWvYNabLY/nEuRjkSewNxOnOLiPs5WQSIoiMQl2Bc8yum96vI1gCrTinHxuNlY+YlgAHUzeAO
gIwlbP/DnHo9F+cUI3MbUSBVkzNttm0ixguu7veEPcihVcRZrP30jOmq0sGZ0ZfPevKBttkspZ8u
Ptr29buVeIKzg1iBaN6Az0PKJfZbHKUWbKz4DpCYDb77rm0aubfTJUwqe5ieRpYCF9Ume5WVbFR+
7eWILwh3IUfXXCEW3LHGjKC/XtvBiQN9KtEl+8rHiW7474j43ddr18Vy949ZLmdpL8WKTngj0lpL
4mVQRBBm4lzh91X0T7Gu1d36dXZqr6pKAyphS2IL/T+kmAVWJK1IJ1C2THpm7IeJblcMR0DUyJiB
aWqK0HtJBfL2mb+zk4di89JS3vB+AAK6SeRssD66rMTD5C1K7W4jxuHYMgokOPhC5eLTLY4JiILi
XigTq8mfhjJwYLI5/92LEFW95pJluskYc8a4SEAL0TH8NbUvuOUAsboU2hUgvVoXmvXk44NsM8Ns
wAwAlzijexMGmg1cBRCbXRtSP4ufBP6rQ/1lqA2KV+TsTzYnuJ7DZAQUzV2k22aZxcTrs35xzzQT
aqAonPunkFlutm5zYzonXisosmEO4hGg7M48i8B23cMiyp2iTDn5xyn/orgYeF1d+x/x6GD9ZL6F
uZPT8bOaUxbmG5HtU9GCVd91+wO8F2uxIV+9Fv3iWbWF9Gl1SLeBujWluIm5WvaTsggbubMF0cLm
mtWowYBATjt6UYec5iNBl5TGyLHXTZ/mob97kpi5ftA3MeGFx0QIs6mWL7kF37pxPF2N9e8BRUEg
vnaYXOeyzLwCg2RS1eevSSc2ozzW+BW5bV4+VeRmj8jM6RA7olAdSdTUluXOLzxDTAd1OPtuE4ik
LX86lcsJjfCKEWJWgodI/M8MpdyWFq+ERnfSQtlBMIVCZ0bYhsMpnyx3hDahXnJgCwcxm/jgg+L1
Y2irbi8XR6B+xMUC/u5n3tQzqZQl1ucxLpab1m84p+nZRwNXW3UucgoQPU0DJexyA0O+pEqYNXMC
7T5GxvztrZHXq3lrm9eUedoEI99TU5flNs5Ibs2CghtolL8cmm95wwTU8/CwLjSbSigiOz282Wlr
sANlznVjgtEiLMamS85JIQ6AAAGADuT97wZnMkXsIChF7Ly1CMDoFWup9ANw7dp/5khccmu8JpB8
ChWdqXrap1Emvubakh97YGjw5y3dEmOjhUEDgaxZ85Ugd6tSUtTy14l9UUKg1Xe4SkqK/VWWYAMg
7LiVmO1zQ9Rioni8UIloqOhXOqD/Zs4mQPOr90iNLMi1tqbdVCP/FM8JhXxvXM9sUHjSM649T5Y8
mF531BNyUO1Vyfsa/JxS8mZaKru3RJPtgevPgKTE/VH96JivZufDxmgJUKYn1dp3gy3TrHJBDf+T
SoVVKwVMc5Z6na/KM1KqZ1dwpRDzb039Zv0YLFHP7bkIfe1O5T0VC6Cu377YHaI99D+L1O3zGvvL
roelCB9YwfPsVO4KIWHQHLH6kVAWYi75/ojvGbnB4IjzGn1k/c+uRiX/1T2lF9GRo+43yOOsMxyP
BsEoOfW4PUD05sMYVRWZ3UNz13iAWcV49BujtaYFZX1+NC30ycYyyEup0oFy5fNZCAUTO+1K+Wn+
80wmDrvKQdFmMa81qemFZwLPWBlWVO9hLQsyyVa/MbFGELKX6TxKIJnSO2vUy7l2bs/iesdzmeQI
UeUxoDszcOWRuFQEXM5x4eqJPGjHuRlrxuSICfMESmI/BJLpP4pPN5WwRy2VCetrk73HgWUxZQxj
e7984GPeTerd8LaCpN9DU/NpHuK8ENcG/43G+lvY5wQEp6sTi8lCWvfEee9TsyYRKPG4/5s1bkrU
Kl9MvgmnQ0XyInC96Hw+Idu2TaD8ahWU8pmtqFX3BXgiWQuvmdWNi1a2ESQUvJamD+/gSM9ain6w
y7WMxHzj+KJyJdjGoTtbEHKtowsFeV7MKaGxfzz+LeFIxTrazDOFKjJ64Ccwl0LzyN1oQ/ABNFOm
bfH306uGSRjFejnGDjHVohxIBtVEH+26lusgmW7WkaXn1mYrA9eQIfCRieHBcLSwT7ANK6CzK3fI
85oRlPpoX4CGgibpjPw5Jyrp1FUjWcftAsn47EHqMkEiP1JDEkHbd8cqw8ZTXa89jSsgOXTp0I+2
U31Dj+F76uHr8169S0HZbRlIWeOxo0FfWqfZ849ZqnfkyjCGOt/oAMfZAcpMZi8ph1IJs7g9aekT
3/kq82fWGVByt04CxUzF5LfacDIWK9LcGbXJwPXim2it/36A2Xdf4REyjR4+rsT4q4Pa3ecgkxpd
Fb4grif2o8cJkrdmkGXW974W+aHL0pHZ6HKyU1ZK/9/ejtg89bRG2CtM3TBFaRaOxg7CmBrCO4ke
N6wZ/j9Od719+btQHcx5iJQ7uA6FZGnXFFR5OzP41ehShH+DeHL3AOVZMHPisJ24VKHXCiuYcN0A
y1RgKQaSBBT7ZWUaHIqozWWwd/h03eSWslFf2Bl45RWdTYmthupFxHkM3/uZLohBi4dL5cgPiYMO
69vDsMJvMHuYdtREuDApir9ERBwaWqZZr69R+tvISl1ONC/4I1Cw9Wtt1uAerhUgqwVWSg+RH76L
aq+C5yVluAf8tENaJ9LSDaEqrtTv8wwBxbI3dna8kqpRxRpxl8gpM0uxOkXaWOvxLamIyx2QABuY
ZN2m4GJF5URNvWZGgRnVloDlaWBdxJQPrY+ghtGS4QPfCNNumMZcOOVbhsCUEs8cGeZN6AWd6pEZ
HKdXZLEK/7dZeAhhOOEy6noxtVKJu7GuPHYl9Ll+BCuMvwLhZcdOs07avjYNT1M+uaCfWqpoH8Lt
WMWgvGbs1ZjbnHPpiGfM2dc3GOFk+hRI9geSyVsOKe00EZmbWeNdxilBhpRt1j2TFdvRh00Yg0yG
uG6qw74K5bWSJjnlqTzpHIgAL9gpm3JgWmQfL1OtCbVP+NRnBEt2TSRs7P8oVm+S2VyoIV8MfowW
I/XkqoKytB5ajF4EAcFseOK3O/vyt4p5HTJrVjAwR6yzc4SrfhUlRZK7RX9oOjY/n0jirE41Z+m8
f26NlNWLiTyvQLk2OqTcddUvr97mv3w1P3KxcHNbxQJGEk3efClkEfcfucYr5rUAzsqCey/rIY3b
Sn4bq4ddXm05qHl0ZYeNx2for4wZ3E/cpiMk1MoU/A+SaLIosUZDGy7PtOaiqPQW6gdczf8ypUFi
iQ5p9AQtJPdY4u/44IURCUnIVgCcOXEmJyGJJzfzrb5PeidVUfHtLqK914GHwdhWRGLojpnXZ8y4
v8eOr4QlH927BldlOJeULwlotp/LENdcc0lnqJAe0PaWoajcw4xwx70lHXEbEfQY/QEaApBDLJqc
qTlgZZhmNQikbpNFczKiaqoD1C6XzdFrAZJpXuXprYGXqrdyp7TbNm2bcGDkOqDe+lxGmRwmpykQ
eJBnp/0oYxc81R5YimHgldZUspzQmTg28UKdAU0BjjQwhe3g0tCWET7MCEKZKPn/NlJz/5OjqOqk
V3UEBbDcnyNA7/JwsJGkgZoRSIRkhNHqhQSIi+o3k8bwVvrSpDggnnKgJysXYrfxGckFWaWs5tI8
ozbQrPfhp2xFlHILdw2xZT710ti1pQ4fSPSNAInTGPXJbviiFyUjYTSDmjl05Kmp7udDyucCzfB2
SZYDEqGAyzMD6oEDVwvD1qEjdTtjc86AsiqpofKjtAqQmnVkuI9pI1rV+rcAhy4e5IT0cckk+fYe
oVlw0IXQ9RD1aZWSKCZ5C9/RhtKOWi5JNQgOTCkUS4v4OOv7oImmhMyxj+7xG7ypIFyOXXkRcC3e
kBIRa2KsIU9Be7ZdleoiuhJRY2cZHOQf5A0Sr2Of7OSRYl/i4CKtam5/yJrVBRfrMJN2vQOGlmEK
4QWCCus0YfHyRMMJtXn/9LoGPxBqgWzFand7VhXA1IeFPJA+WLsbrNISLbKju9OR8VXoon6oO5hV
OhWVpmjhtTnWci+xiipfmPIzRT72D9Xnm4ulo5VIC9mY2+1+Wfw7MDn3NunJp+XCQI3CX0NazbnR
tyFirfrxQGprAz00ex+rchPoHgSmIWUBmmWX2BnlgQpR4Og8a3dFKNwFLTS7jiCZJyXrqaxDSubt
azLqk/vVhF/Mi46s/CZAFMNKEVyjNHQWeLiC9486dmAVmFTi67XIXn4vyKXh7LjBxlSNKtpatnD9
eDr4JtPdwlWKxvIlasgswfSuFDV1veSKkI5DCjIpKpI3uhFu7LsTA7gP5b8iC+oSCmJvW2Othwut
fUeco2qrFqQB2YR25riLV6BNc5DvyrDt5XyQXZL9YX2jkRO8c8I+ExGesGy3WQsVhhCgPecZlJTO
m20S2wLji2bzwHHOZazH6LV0BH8qaqWlLH4LmzCWyojR7VhXYfq0xx50Jrx0ny09yyRXsAEMdbeB
IAB/O3YIzhv09TF7gvLiJpMAN/aNRhgBbUxoTmaKa0MBxiwWTEZeod04p75y5SWXACzQHGbfdqHP
vhlA5RzXKMtwZ0m7sDp/EE3lSC+dFkeyq8Bni0jUT4NcH6Rd1OW6GsgJ8A2CKaAXVhlhg2IgPoMB
9ylLCYXnqyrTqZDghDfreyHNmu5zajhhTw7MEJEjBW8C0oeRxPjxdEj9nezwJ9lN7thA/rRiwRwL
8nO9CcbSy/NEylZDCPuEG53TZBkEVDaXgzwRNgyvDEwundKQ3iNoyZvFgQrbgrvVQZLaRhLZbn2M
nSkkMid7bxkVzkdzO6ZD4r4dolRXLFGKGChTmBYs5kBK/jZqB9U2V1OSxFDXJOOyksvsc+Vm3tQ/
oC4BH8kv7GrqPDfH+t2tO2uECT5Sk259EXwpqF8FDafrJfoPzXuvgxh/wLTG60vQJMlm7FI4WaTc
2u4lxW0XD+yGquQmmEmmJyiDNl/O0Ak0IUwfGzw9kdi91jxlJvYGknlO2uufL6v8zEgPmNsc1YG/
IvPAE7KEd3AC6Zez3QcktrSQr011kzRILUoDTSpEF7DdpmK05qy+RRZOjcLvzzvzZysVEHGMC7/W
Zy5szi8DgWYC3zA4bkoZ1SWmg7DK6Ym/5oW8Lzh3m3PuIZCMLZTvICiS59TVa3MDoeD1LV1GFRFO
8I79JQZ6i3XtzwArTA0fLoAz52fS/jbPcsjBg33AT5OeZnbAYG5B3qtI6MyoRmJWzM2wmkTKmtQp
1r50zmSCT9Cwxth3rWpn3kUH86CWUonlzBsJDpbBe/MV859/U6qg/n26NQaAQjsaW1lpG5qI40jh
PGRKxiyV1xW8ZNqXbJUmLy/A+WOE1TETZb13PB0BUObiPMoWuSods2jJfixGgEL0c79KX07UWAWq
6UJHOrc260n+q9s4zXt6lt/Jtl1MNF5Lta6OKO9BQhB/grqGDo4HFgPFlGOauc2ZNHp9511tW5sB
MlU4nMNoToRcONz472Sh+BtG2sJxBkeuG8eunf8pqYlM74uU5A7mGM0klOuiiaVeRVzvUZtH2+ku
5U+juhBPrLzC/1IlvdbSUQ8EhZNAJU7ADkKKRJ8Y+Y65PQrDjQddB7munxlQV6BSaD0k5BWVg7Dq
L86IBP3vd1ZgZ3c5Y2TNprucM8JW8jiDDbJwxOKoEq5D4AMvNfkq9WG74o7qInZQafh2bRe+Q8Rl
O5DUosku2NeT24Czi4vHVKb5UvCL960ss3Vci6kOCJPV1AkQIP/qQdgUFj3mrU0uRg7Pa19dwopi
S+b3xpoftnRuRsS1YiAMnAZYTJggPibIEKxNMdcZWRtzb7tTDqBfywMS9zCCPJSkxw57pC8TwQaL
3aaQDUw+qYvIv4/lBhmrHPN3O2s2vKzrQQs4HRAVQeehXI4c+r+2eClXI32GXN02lyHJ321eqlG8
ohGWjtxTq001UP5hclakFf/bDS0Nq6hdaizruiK4xiJy51TApz6vWZ3WQshOOwxf1CTQrPCx2E8v
cEE9RDTK4hdLH2YQf+qGmd9tL3wq761KQqnd30OV6fxXZ7eYi4h4b/riOpiYpOV3kEGJg3ukDJ0l
DatoRDHHcls6tnCrXwGu1bDt7QbblFxAac31+Aqb8RXi0vHlBR6JCX05KYTdCuoyROjOTYc624Fi
oGBMgrNsOYi9vc7Xmb5xPOyteHo3MxljGL+cM+64HeVYVyVqPUY2a+6mAH/lYhr8IdlmuV3Itpfs
0hb6oVxyd/9l4x+HCSvw3M/gYwqeH4hm38F8nshbpjHpevtAbgd032/8ZZiaVNWcfm89bFfuImbg
gyK53u3fGa2O8KqrCqvdRsoaje4u7knlYHYFXpBm09QabISrjdU3vf70fzqvwtQGNiUQ5FcMXJyv
7OsU33Soh0vUR78fQoBT+fIs61SREKYKepb9Ui13SWXveesrDFLFur+4B+Gb3MJlEZxEROU6FQpE
pyBIrotB9J1Bl3KRhZWQ7rwJDblKUINW3dqTQNA2sTg3GzU89/gqEpShpE9hXTQFTAy6q0b1/+8c
htciGr2i0InZZ7u8sElsAjttXc3AMEJ7xdnaBFc5+OzmhfrqLjmZVI9BG9nwI+5xNgp+6vNLBiN2
fL1LorMBp8G0qj31fQpLbgSoKM4DzBP7yz2HxqbeVV3NTcnfNn46/gGCcwZW69oPlztRoZZjVgWW
mHkJP/zeMVTloJt/ZHTiiKm44b5tKMksZ2bwyhPGjQLvII7QjhFIyo2OqB5OZdQjkEot/YqfXa4w
oxsyAHrCMwRk3iMu7m1UOGoKvOnspbFo81mDE7Ihd2cQEzJvLri9bifLXxcDy1XLpIYspIpjMUZe
41PSgvbJuUNspmVAVSi5iyc67Eo5/RneBsHOwshRr4nFvkQ7CUcS5/Tsp1RVJwLdtcD3Abx4uBgw
7Mjxuc5sCfo6xeGAEv760zMGrR8lJWfFUN/i518e1dxzre83XjEAFT0rp7NkD2Nbtl8GIkG4B87A
uZmWZJQPEMMcwJO7tQniXHag9J9+2trh602igxmQeBuyymxNlJy+JA5VnLiA6LFueDk4YN6d3R4j
XmyNjNb+y44fnhG5H8fBz1mHp8nFZx9+GAFXnjbqaoKhd8ETvEXYnNt/47rR36FzKBn93OnCSYR4
fTf960UUvkPWLDTHdRxBgN8p0+TW3t428/62y7fesUC0LEHIrrx14zGWt5M65dks5aj5aZVfiVr+
YNu9oS04BTSl70lX9JPwwdOAV0YnYHtd7cCIbtkHq1uhHSumsgCHa5KDKtI/SrOXxlAUwd9OLuIj
mZnqDQYEwcdH1wdzk4pGrDMFKinX55srP7/O8++zusVkydCiqtdr2U1KPhbG+O6lfIPUFh5+0Gks
lirREIao+wrIqLlI5/3Y/KEWPgBBLOnMF/p+AckyKv3TL8GNQ5UiEAbdTbozE5cgDq+hSQLQoWMF
vOE5MtVdVluFyV7anKn5bppG2QMdBPBoTpuK/INx2ukpO2D6ZaNWounD/jRvaORK8sSniLdMhwvF
pJ0LfeYliHn1MQGKsNOup7OJbK0OjTrAn67ekpeIU174tmY0tHf/m/LDedKrT9qmEotqbRSufrLY
YzSs6xpnD56//9NUf3vdID84JSLVZaS/JOMJ20cb9mDU50ZxXtHFXHCmpCjn7HX9oCLe1XFDeMmR
GgnJyz44kXw85Q7SQ8HdrzloQFT335FPCNKhvML2vq1uuv3prdXb9Zw7RsKOAtA3yT1hk8RvtsaO
eply7niUoas/bP70rntskza0foDm6iXOjheE3FU8s3NknO6uuTPiTq42+NOFFszoYOYp48EcFeiS
V4PB/IUBjl31wRvUOR3EDYsy0klk8aVg2VrV4s001olkRvcjdAMk3GpkkXh5H6+eqPM91dnSMxhb
maSTlHcvO6PG4OijcFzeL0GYg8TLqjcwEmz3GZq3RV2ukkgJi276dWWKD0zRtp3Zz3MA1fRZdxxv
tY7fK1y1cd7t8nmD+IXmuPT9BoYaQiSI6XAUTWXGvRphIhLhagds8SuM1rO1oWmfMDA2q7f5x8rZ
cpz1rbdkU5nEG3ztILBxiXduXb+JeJhegYjPCy4jAKy1tay8K9DvoTlMQdlEdifouk9EJ737xk27
7XVuuLiInAblWJOEhMB3XSUVMdpU4NzKojh3nNEXzYrgFiz9CKxQTKGiMOwVF7hUO4nD+c+FVeB+
pdhxI9KD7q7idU/LLg+dYukwO5ptABz8aXg2ygDPcZ7J8IXV0CK6khX3QeUC7fMeJUomATTMGiwi
I+FNLBMdClttK2uESvXNz6zcNvfDkyfst1aVqLx7ZE+h9bUtDLRS17y9Rn0w6Y9Ko7t5ES7Kf9/p
dG1Ji4aHuSkFE2yZvXp1EpDzNM40wbQcbxyk7tSsNbnOn7cmwsAac1KLdYUvcK6AEDdYeR2SJa2L
IYvNGeZNDq+VlvjXAwbST/PoQ6TleIpBj6OY0OgpFD3umZAOTVcr4z40Bgd7qeLvTK0jMIUgliOu
PCkE52sl+ZJHXCxwgx0krQPPhl/eoCY/4R+f6UTEzNiCVnHYqHlng4RT51Tm6J2dZzQN5SVi8DXs
/+DS/+jfMgWPsxz+zqJmWGjxGSNopDeLsrN8/KB0tBKH5tzy96a4PXjJv4smZZXKgbqAVyFHUQsK
HHvSoXwBXyQYY/Mu+ujppHn3xYrIrX6F1VFUS27gl9hZQfSc3ZFJ7/G10faosfX3ffWk8+pgQYhT
LThyTvssHH55kP60jjZphQiSHQoApZUUOVuu4bJv+gdujGqbasi7wyVCV6XiAYZKC/bX5PpgdH5r
frU4dim7m+G5j42KIBBzZdvUgCBefpMQYzC24XPWZybqoIFbQ8n/pMAWwSmsLiUP3uAJsPWJd10U
2EIruwsiHq7v5w2eiGlZc8snyjp3pZPC0kfXUI3u34hccBN1WKeAxvD8kKTKoPiIRG7VM4hbF/pP
uBVrkbJI/Xum4i9ROroXBp5vtxmSStEeZcLqNe5+9oy9PoCPrxjCz8gMHi8YKS6YT0YdH3xLNk9v
6ZHuXRQZCtwazoKzp+XkxPTy0ZS5qKWBj62x+OwOrzBc9YqDLiJW8tB/tmki+IoR7YGWLy1dDZi/
aAbqYPLNRwHvDPV5sDAyBT+Rm2ucsvYjURuUE2YiK95i6wKkrTRFKvxWAh6229sMFyK8kcWl+JTD
FexvjtFQl2XbUzFFQQ6r7y6GpfbTcLyUYiMw6/1XJ7tvg40O8Q5gike+5yEeOr8S2HesQXqDjoQX
pyq2cuC3/iu0DtcDG8dUhpTHelkT07MqjmDG/KCeYIhXqqshFUMubjpFS1gYibK1xN3RQAfw79L0
eqy60kZzwVTM+8jxMo2gfyvMm3IfwI+OomI5rWYf3bHMyfqFKGE4v+/XWHMw+vdL2wU+TVqZhtgN
P1WqQ0bSPriWKAsMOT7/EswJwTvJJnTmGZB1T/ckUhrpHPb1j3/0Lrj49cmjGIMo54FvfaWRvpLK
cXXeKxIMAtnYGzvXmXNfZfIbwvsoCCHe2Aij8ukHCISE0I4PmOPHgfbEZoz92OLBpUB+b/h5Meo5
yzXxUt8A3SmioGCwdVs0ilypHX1B7nz1+TQCv2Pn4PqhfIXRzuKZiS26652mwwio9EVN1qBQopqu
nT0Ob1ee4ryA/LBu/1sOyIhtZHdzlk9tJte6gPwOne0UhB7OjJnsKgpUpDDTYZDCXasS3zHryOz1
yKVPz6papcIjsrkQnnimC6Zn4tbCniTb1Eceju6Ig6/ENuwLx3U2JBbLHyu0W8mYQyBfJ6BDbvaI
O38oTl3QWKjnvnTtMAURKrQc3kq+x3MQMm6M8g0XBU3BZvkljGq4gPjXQiT4fEqd3aYXRYmZ9uE/
plyA5PCHSIRi8UL2MJw+0d1SqZ6aVnzQ6gMur0UCCuBttZgezb99XWTS0jvWFeYMYwEj1mmUYUb/
7h8ktY0SETkDe+Qfeb/DAs6Rp7jKb1mQGLH9HYlz3Tc+hOulcDZ/9ECLHIPmBubBYXe14w2Blggf
8B/oMlzt3ItmE2/LnsDarLR2EdsCcS+ZCuLfGagOdChw/QP9K2A74Pi8n9bJjeY61t4qAUYeU3rF
3alvYOg1TFMwvAeyjK9Jqzam9yesZLTctQcmlA8It50fg976Gb8bqZ3cQVYvGNFSNpiKVMISCQex
5Vp/Gbz626qeY2gbA54NAPEAwhyqqv/v+SAWbmh9oFMvyzZ6EXz8D2oLY1bNNel8kWBMiogDm8Qj
lcA13rMXZy/8cz2qw53aQX2gaABm1NsqQ1VSCCCTS6sjReA8oqVKCANqROYYoHUzoklojcWGryGT
EY0JymrHxsMaUohIw3Vv1KedrtsklfT7lKr5hr0BaamxdE7Xjuk4R5pUBviIwNCprJpGBho4F6eO
Rrxues+iawZ7ZqfFKBmf1JR+dNvGVFu0QS7dNXKD1OdiqZkK3BPktvt3kvA+oqSWG7BI5QC2t1NS
qNc1w1nvf1glrqDINplO7Cozu7oavtNmPjhOu880Rzg4qockW0JS8uLVnOcU3+gRF8nHj7RCDQWM
0s+UXFzLm0SkDJSb6R8A6OJiBJPsa0VSFSgwTVuPpPr1hMDCrG3Ohzgo9awFP6yR/ZwePW85Y8ND
LA9b7eKnagve77Xdug+uMep6jZPNhWWHzVHPS7LWSo/50GePEAISFg0Be7BJr07ZKycM7VcJV93o
xn9AV+I2zePDO4SifrXzXiMnoeDrUhpB35C2q1a4eGMg2/mOVoFljyLtSVxucjzC+yVNv6gtlk0E
ycn9+tsu6cw75U79ganR01IItfQPlJs3e9SL9OezFs0Ze8k6x0z1u9VaKqqWY9eVnQPMZnh9/let
JA9F5uahPlpM2ol7ak3nzfMJURwj/Rfu8bogrHF0SpxVcGTD7Ww09UDm+1bbemKnxEi1GzgUirV/
qfRmF6IGYBu6A3Thhgfabvkm7jBtxuqbIfDxKbZmr+eT9cmUKW+8D1T7Y3LzD8gKn/5tQLsqG8lk
DFGdtB9dAnWeOrp0/pYW1DLyWothz2Et7P4fM9Sm11JdOH/8bzm+FdeL75XwhCb1UvyAIPAMPVi1
mILjsk7p0m7hjANWmrfQgCpEKL+vufmJzzUla8r9B+DCpTdH7UbE0aGJ4LMvYWIPVsYrObpKxuk0
ixkMOZULLyy0kN1ag72pF5KHEcEEAf1PJGr1W1YiIas45V5cmmkJuJ9KlaZHAKKbvOcf1dNSr+47
zK5yb05B6kluWOevwqd6xWahuKQIazx30OfubWgbGCEtucoP+geEXzPgutQO/epJ5ai23TbI1fKX
H9VnQyJux/eNpvB+DVI8SGk9cd5yAlGtwT9zP0YqA2SObIBkjfIiXv2ZFfkmoRoF9MTUBaXwG1BY
04OBpoxTyrtMi6O8W790HL7DxBdbB+idLIliuFGQy50CPKf0F+4uhk26msPRAOU/3faZTD5GlHee
03DsLnKLURruw0qebmMKrM3M7TFtiy0ISljDyQUhX659RUGSN1epcCJDmUxw6gu1Ng6KbICbc3O/
Pd3m3UNxWvzxeUEfQrqnl5KwDKD2htIVSeJr14qItxxJqwX2xZSYgP7/FzPq8Ak6kOyJf40gKJvQ
RLSL0734VPGnYkMEb70fkqK0/P0f84LutIFEVAs0F2DxHlAJBVawPOxMskmAdgJrWEgGKn5Wb62w
Z7EeSqsvU/5JdihrW08mJYTDYNFnPLqNPKH3ALpOg3lCTG2+2/41q33lkjgv6CBwhA8eLTNwGpLU
j1wKhuWmAnAKbhQc0iaouSWkEUwTIjlMF32kQnpdv0pknNzl1Y5GBHTborrVZbzHL9sJfF08lmU5
PkQfPZ91EO0JDrRauR7wi2jOyn7I5tHjJ2GSzgAdbCKrsZ+ia1qGAq+07K0i8xzYYcvQwKDY6u0K
4X8+reT/RT0dgL3mE4EZtDWjI3mGgBiNcjjBmcDWTsjiWJZ+OWs6XexH6AfUbN8JaN2jf3reSo59
GZIKsVbDFBXEzqSvTU+HYUI4v9D4DztaEWck46n73aJMTHdrLN5ZUo2R38tCg66XAD1ls2YNhUA3
7wI4+TpAjtWMKUKSFbyVwbMvIvGmRonjlgA9sk2hTlgBvoeHWKy492pDgTHtUiQ7wMtXBSO6LGhY
9JMMrUwQf1Ej/5m6iMleVHsVR1ehPBoAn/9AO238ljKZ6RZ/xP54FGl+yDJrUe918fHKFFq/j1EP
RP4x2T+P/IRdhyQig+457dAPe3K962JC/WbT2y187Xm/uAaRuB2ysl7NBanM+O4XjhFoIzWYzsQN
AI3mPbCeC3E9ltYOWhCJQmNHNUSRGMF6NwgNvuQ+v/INXVK33VN0TQw22Ocb+Hpp8RwC16i1CpLM
V6SRIluOIawWeQPuCkbGplXaqInXOMz6FizvlYmb+hn6d7CtWkUOuqqMIbiZHUCvp4VFihkz6rqd
D5A58gCVb8Cqjk7FWFwtT6+YaEeSDmgxdYb+Hd9QBhUU+G4zvQjrgLWhL84CR3mClImQEhKdJNre
Sx49X+dEhs3+hBDg/ePL9MLy9AIrPW8STN+c9SDkrAaBhjvswfDe//0ODU1dVcUKhKtkdasfgbYs
/oVdmdyDY2SKQEaNshZU8gm7cvBj4G/QnmYlSKjdAX4C1Vam8tj3JfBgNKqOs2IPM6A59s1J/8OW
aDQ5pU5QC6Wty2oIYQpaTB0AxyhBeZS0Fwd+s79jj4T7Au/seXxczEeoTRjeFTUVEeMSHLAKanCP
IhUmoBjUaDfW+d36tm/Ilg5SUbpezZxgMcD/PovMa1TmgKY5oZ1ozgotLawAABlsupoVFoDm6/eg
fAzN7dI1Ooyb7B4w8X1F5Oj/idm1TedW9tMjVzKMANA8xzRg9taXyv6U98AqY4cqZBnLzNgp49aD
sRUbdeth/eeqBy/0Ksc3gRM4b79yWP6sZc1E0/I6QxhMVgTRqeBrXxf1YSJ4nScIr6V09C5thSUu
dQQH/jsUGxVwqC2fvSeys9Vf6C7NS+37iC6a3CA20kSaDmSSzPsRy2o2fZ1lcoh4J3jsFfMpfH3O
kD7b7j1RrQhfJMaWTk6LDztU4rU/hOCx6LddQ3wbfzaDv2nU8H8eNMZ3ISR+fIHXn0xCQWc/ITbN
VqdgBKh42aEBkgKz1SKpNem7fZvrtDBqiUgBiMbXDY5F4KAFEynZR6QaBb4n5u0+bbYi91bl2Y/O
5xTJtI6kwzlvWHAWhIckYm6tCSNyTZTMDJ73KBSHR8HwiasXxLJWKBQP+1Tspd3hLFUnaXAiPvXZ
ehDt8Xaeppya1EeYdsTYaJokzymLDhaTo/Z5fgg3C9S6OLOHxi9P2ULWI80t6EheW8Z7SqxyU1IK
xlUmONgcp2dHR54IBiTReJgfTLbpGX8fGL2zZxLVq9iSm+f4A/zQXgTKCLbL3qm/HbWoMr7AOeLE
8L35w9089mv+Yt01dQwF3p+wSOGrXqmAQpwF0yNmWd1lEV4j6PBgP2benv9k0yPhFWxPBxNzFqPy
Yh3YJxc58FkWzQsb3/AfK9qFsPai/T383/urT4PiM81XWJFb03P+Lmfkiu0b3543JFo94Ed+k+Ss
XEFl5gnn0mrirP5/S22q2Yvje42SUGakopD28YCSt1k9k7Y7sR7YtJSekymJTK5CSG3KsHxutOQP
CHlDPPaRvlHFUX9TDXi5uDobepuM6ePCs9ryYFsn/7ONI64ixK5rii30tqmVFWHYJqi3DSCcOkBb
GEbMBQiQY69miUTG8+7sXyQaZUOjG6qUyOlq3PGeWgFIkNgNk5JvT1F24iPgJr8toS/ViJhhgy27
4lR3lm2spocBOZpJjHu/Vz4Ki8nwjfmMWd6kaUgiBY/wgO7tispJ/VuYgMGWGKLU7oSaXno1MINk
aosh9FKfnG4xRcmwRnyglMGx1b9I7PUi2iP/rbYslYD7N4QvYeUg8PaZMSfJqOKpYJOYUoW+UZDS
diKW0obzAP4Bl5gN24h1NVihczPLEvsUwrSYpCLqNOnwdQyaxEr9PetUKJPfwJZ+IquY68HZIzg0
rQT8/QwvLtdEeHFnsiVeWXI1RygigC4xuoGrgbq89qWEtx8gx8rJ1ymF7amV6jtmPZK6bN3bxx7d
V7XzFgVNa5BClA7JcK3BxNWsWivNT2pK4EMNuwqDVg2FQAUbMy9gBytst9CPvJOhdT+Ue5ZZSdCI
1i7oW62xe+deXNfwjJcfTLuB+JDaX+1oI1c8xSxhEl8bVDKV/8tpUPwOL0C/DrawRy1xO/MwAkSX
2q+Inj7Yrb6f9Kw99McP9xjpc0UM/dHD+L6N+utirEP3ncypNYS0b4idUSpEr5gEQ7LzoUmtQRRu
i71N/JQdmkYA+nE5kEUViRhHSiW5vC2ssyHrDHH2tjjI2mS3jG1MLA32MgEhzdha26CHpeRa+eiz
Cz765bFEypGNGoZtsAyn8EtmEHRtIokG16xi0R3LoQCNYCo3gGJqvatlrrlk8c52rLF7ifLn+nxI
hl6mWqtDT6wFou6ZWxKdU4t/JyZKAurz3NLDSc+U/7o1JHp4IDL3NsqvEzm2aWQa9T+AabhqSGpM
PlYRieNEYO/IJAdxMdOfaJruTtC9UcImOYEsEO3yKk1Vq8tlo14/whZvXxW+QcctWPaaFdEPZWNE
yK7GivokrbDC/cAV4ehpZOYp4wN2CBwaPv4baxc+SwvO+IpPxu21KxYFSkxQHFe7/qaS5mf5fpZn
XZHgPo7O602rpr38Vsx4NgU3lnjXFs/DEgbA8AQyYeJUFJT1senOYlXEx/Wi28VCt1k+j/4dk+K8
Se8Yp9OyrRyopP9Tbv5tp87eyGXtTjQ2VvxwC/H5RhVg/vyEy7eoFI6w9FGPnYQ9HT/gCRTi+axR
bRxF8dZYxemnIxQSClw+qkqWR0EhVQ6W6GHe9v29WSNEuV4hVvipbslD27HXAy1Xk6dne9yEaG8V
IO/7rC/Th+lyCXLMeoXnk1VYGWJLABhS1us9KZPtvUXgK0ciUvk2BW6ceGjlsS+KGbj5SoAIr6od
tx/TkoxNwV9Ey22UMN3gIQlnKDGYUiDfSrRSZzVg1lOmDya1qDQM0sD9ZyX2RHm1bBuGTOg+0uN7
t0P/zdjLIh3EevWJdigGvaFt2N6buoM9hAuaCbNkGt54wKxxDYOPNhRJmg0gcmjGg40QTSlcVdwI
SXlMfHbr35kVi3wg84IfFhDIrWpe9QdIf7uEVoFupFjYrsQqf4mYWSYQ6ItWtrMmTqXV+43xr0l0
fQtUR5Oi511zXDlaseHmbO81jx3cZK1r028ok7eI7y/AjWMTMF0fZLs0XjRhHyxhUazqg1gY5cHh
dUajWn8acMD54uDuD/UBU69X4GJjY4FicZ7AgD/V9PmRoPjGT585wxIBAy2p6xjQtehSPgMqjpXP
7JUa0LKJSTBLrQpmnHUum1my/EUPtzZ/2R1xs7fm8Bf4Dpz9QafLXgj1HurYAby4WD7U8IZg+BLg
mo3FWDFBBnMaFoo9rS+cl0sbNVqPNo16RyqVwn4NaP/XwTWEpLlswE5f6V1nQ3mP0SgbuoryfO/L
LEzU4pvN9LByiYuPKx8ydE/x1wxJIkQUIzT4dTHPcdBa+x+vj+wVsPUs0Ay7jIKcjnem0Wl/aWvp
skfIVwQ6dOj/jW5yDkvVsoigsrNDEZGDSKy2LHZbdIEOe3zCe3WzI4LZC6RApp2le6EMEvwcckW/
xA5rFFgdR1ts473zwDLy4wiRbEXMr5Zg+6jd2jFvbVxUhq2xu/RNr8Uzh7rPqt3gv1drhXub/tpt
gG+vT/rOyy6B3iaeZ2qaXJUVw7L6BlHPw4XtZezwAKg8c3puWfs/8N06EANSQOCLMHQNCjCCRkU+
9bcdwVKQdkC+Os4ZoqFjCKnnrv32hEVCJ9JD/Lc4LMWQtyCbR0fv5TbS86d+o0q5x+BqrdpInWCq
7GAcdEIkFzKpvAm4A4e9/n33ZHeYyHlE07yyTacc8zkj2fzdYmx3aFyzO30DVgV0qhYKk9Q3+Slu
ylT8yZ4i4tZP3ZAE5EnXrAJtv0AzutDoZ7p8l4WSVRyQMaepPRn+2rApd2Vt9TqHRyHSpRniFNmR
eguHuQ0qt5o+pm3LCeL5s8TPZjWVNVgLvP54Y/iellqIAvF9Ddoi5JaiKivBeLW2dTAqRCl8Q5cv
RN1XdzDpLy+W5EESV66/+FiBBKhSZPNDbMyQkhncRCYD7+s3rAKPsJ9NmGjaYR6wVHGANuAk0M3C
S4XCcs/iDjkbneyBV47Az7vqUlVfsLmacJ/a22BAPuCK9t+9T6aYTwNnitlQcKvh3c/KS6fbObPo
OsVLfzKWYYmQiq19i2cEikh1u94KseWiqrLrgD/H7nmfH2K1LpZIzPCW2rddc3mE2VXkCa5ejtAT
Pfxegxij6DrSXAtbzLc2VXOvimSf2GHtMVmA7W10FVCYB7CsajnLm+D4lp8guvF7bmYLiaXl8cOQ
aF/XiqSEWS2tJNEoIxew/nUkdfZgkoiggxi/IKSAoymkz5kcl0vZOBQ8Tpoz4s1j9wkVJ1h8cmLY
Bg9DBm3+Jl5LMaxmeSAAmPGhrEU/huFWgC/6TdksMYq5klp6CLDiQj0ABsI9E5j1evbsoKb30B+a
2d6VEJf7Tkjd4/H/7I3ElPmBpVPW6yZfrmwS+bK5grNhZ+MFr8qUXIkwOqv9xUKfijDEmqEFqpm+
6Nn83nVsRpjtQx2TmUW5bB9ecN+avTfW0jlavHELMs+UlH+QMhuo1/2eVpXWLW2i7IE5cMNwNBR2
1XXWFpGnMC36ZqJysjyBgcmSHMDYljxhFjYnoJx1mGlpnmi/8hvl71SZ7YDzbmBY2S1cU+PHRn8h
bjB2G4c4xyfywSoJwitaWNZs2tWlo/yc9m3lBh/pkm3tjcti6t/2QH/JUJmPl9otGNlys0CWzqnj
CmDURm9ER3+/k4r2pmKGgWRN28a2rNZUxs9QIS4nyQ13zKpLj9ZsRA/FrTSTPPc3olveVzduhvKl
OdQz3BptQ6NymwP7jJmcrwccYsxJDOM7qLVSWOnKuaM+Wk56OIiJ15j/LCSUJBKkxSuwpeHp1RlG
mxXmylob9xs/6e1vKknDma2Wtuhh8hWwKmBAzaS7H38zhu0ITdxvl+tFpAKBKEVG9F6R7IsA41vI
ex7xlsM6QOOw4bIZZ6iUYYQlSvl7i2ZYnhwUWJFBZPcen163Iqz5Tfxa8GK7ck+N2yW/k4pgomGB
BUqe2NeNB4gYHX7/aSzE6/1JOZYi+QNkdG2pmiqG1AjByP6IOcVSRQ7EojBcGNZMWHfOmmXZC8Qt
YwwtSSPzH4wy0XAX82V1W/otaZNpZ3kSZeJGwzBTzDV4eS8V3s1+MTVvo53LPl4m7luOKiRDbylF
cURc68TjoydX2A3DZIfNadHigZNdxLk2e7s7bOA9C9UMrNpDZQBPK/p6u0koriv5YePeXQt5IIO5
wdX744mfqIpCfbP5pFGCelx+AkHwFLGySEdnr6D7LUbaq1wTd6dhO8XOJJ1oos5FU5JFpzQ2mFdx
HsU6TVaZBdBUZHvZLs8CBim7zz7/3XSEsB8g3SEwgUqwjdOy7rgJBvQcg7yVeofGicDl09P/xIA3
g2rKZczh5rRQT4s9Y04LgM9OmdY1BNZNaMiy0svtUSpUl6lhBawJhRFMwJs3LGMc9lWkVrvdaHF/
ivH6Z00xQJ2QsOsgyhNmlTzifLnLPPZDiBuHF0YyPXZVubbOvpsOsAsiFDrENSFY0EEodihyK8Jd
coy4JEkVKB0u2Y1n/t/NWBASFTD+YJHKd+iaCi+5APin8ehowWExRwb5Zub/tVw2BrRWC0mqiZQ3
Qw6ajgLRjSg2tO5Sg5P35+hrRykElMv4zUBqOP0RRI8oRhIc1YzmEj5ZLlEFR8KL2X+1bQaW7+8T
Qp8jqRu6ilQih9ITS/YtY4Z6PT0g1eW/Olzc5yO9nl/sw0mf+qfgqtEcYApz35Funkeigszdj+mH
cLKnknnalmDagbeQVyULV2TVEqAkzRk3cykOYQViA+zPAZj7GdDwzql9oRg2YHPbJDn1xPKz4+xh
Srb3eMH47Qxqpu9hCVk3hXRZrtdMjJC1IWN/vR2qw3F9DIEoJUppluhTStsEp+0Uw6KwNZmg8MkZ
+jCq4IAhMnRdk1f39tHpt0Tx0F4gwsqj+cXJNOXZ+l4g8n1dVm2SLvlgD9ADqozy/LeSGQ/oeFQ4
4JNF/3on7G7SSBbk5fHELJosj/QlZirJsZCBtGX5jr5BboP2eggX7+2KinEIEKzx0fQkBRrxgnEX
mQEHY4BXUG9S0npXQ19iFe4PQpoOqPc1HlDmgakVbKi+FkRe22tDS8JWmTjCweiJld7/0DN1TZBt
LAvroEARjZRcrVIjOGBL/BltFKLZJ8uUwOD3zVKCZXoMXsNhlEAxtsujrRVEsR5yt3EBzI2s1604
S9rkdk6RRqoNaUznOMY1BW/6HEJOSQyXxqavg5myCGgRstdCCdtF1Nzehhzt5kgQPuiP756/1Lm2
Wn3GYdYOrOVelrD5AN0uqGtbIXqCKCCSjXYKtHxeGCH7/ujclklpCeHBhY436OG/QS9dzjiA3r6R
WqZ38DnBljh25JY+flK5Eh+PiClqduhOO3h4ggWnIWuoSVfz6w7PSd+qFfBCtaTJzmAqlXawNBbV
eo3srLBip5zuQSOojofF1Lcrn9LkJiFcOu+oUVK68xpVaQuQ5WNm2eeWq9L4wSIoKJPgLYzanil0
WQhOeUHi6rO/Hqb2c2MC2sYSqo1Wy0RjVqOVi9sm0GqENPVXDURdsJWkmgWGSGM5vZp6NSX3WJVt
s4fjZzQKfLrn/KvZ4zHbKHZxWhxTj9P7/jTZhAZAi2kdHMHcwWkuUMnOBf38U29PA6q+DvgulXTi
oP8PC0Z+KtCIM3Msisd2O5SKNvsTzGNtDJaVwIdGXQV8fVEC+0tiQfjMufNR0MApnfJSgV1bRKqB
A0aooA8oVAZUwiinMu2UZhWWb+aVD8HUJLmhqMPxGgb/EeQ7JI6dGNgn+I7XJ82CO2O84DF3MJp5
LklKWnMJ3pFXtQkeFEcMglrQTs2hnv9MUhR/Cx7rFp17NEEMn172eI9S4TsEUyip+npOvSuIvuPW
yQFx+0wGYfAkU36w7k8XqvnIT4Nb9rxRTig347nZQEa8IJ5IQe39VI5sYb4Lzbqk6KPvFpeIvDIC
9vNOqdN91lFEBF27gqhUc7SnJq3ZH/wS0uugYvWxA5iawCbCiRY2P2YxdAxsiUrEYgV3VdYTW0BW
ebrrNA5jItOv55nspR2Av3QIb4ZdWqrtbQbJKDqP6mjD7sYMWyeoMg+ShKtIAz488BQzAsTGJrvc
l1vo1N4+LsTWr4v9aRB8ojTgueUs5VfLJspEyx86ukD2SYKLf/+MQMXeP2wWvmPoJHV2cfSgoqkT
RccJnlhOaWvvMf7xMx2UlCplbuU5hruCCwtWlVV42MVAvWg/y8kIVJYmEAH7rIy5O0frPucyu5gk
VRU514n6Q8iKYf/QDFHgBOVtRyGIUMhfprl4qf5jTiv3f3iCZN31jj1ieo7r49DAwAGQE6zatlbA
SXx4x/wreOuvvtseszvN5lJN1sSRER37QnCsGFqDXlXKfGG1S9ApX+xHcWFIt/Ft+ZJCL/iXwM4y
s7kNtYf9e7wJI8cHfMGpOVXCEcK/Rx/pFiS7eLqnrW8eKi111pmlkcyJ1aG/TcSy8B6er7m/rg1K
GTxtKJPeCpVepxi7otX6qRc6VRoF0aBsE2VXJjP/48rjud/GaYQ2FbEqbD46sHcmjdPjfFILNdma
wTHfH1MoIdn24s1K3YQON1qBbGrAbTsiRz4qiYIC2+S+KOczajpeJlEAjCJrijMIVg+z2DmZtJsh
0rUcsg1XkQSUFG4p4j9ukl6we6HMCfpwwEhFlmVSc3U7z0UZEHHTGj/BvJdoq6vLaeYgXxZL5JU9
/+msXoThhi50IfA0foNpHS/9c06mZsu5zyeSzBwgmel4CFPuImwamYCkJ0+PM1ZSRHEeBq6SkzVT
s0T1JdUjyMXtmWWC1ZyFKlVHCEwNbYgX4is1zuyuIOEYom1XJWWZwkiCu9YnpLhzbLeaXfkoNWKn
n0+STIfe2wpIpA6xdKmNEw6eRE4aXYt3Qd/2LpjdtTR6vggO96lWgdZQcEyxiBZtdWhFTIpGFvfq
L6YxMV2LwLhjNwvMZIzhoOYsMl1+7ohUen0iocMstOC/Zgd7vPGbUFeg+MdzppDNIfaHGEsq/gNb
LzET7b4WThEF6y9EZEp72GvkVowHsyfcWksSVUuV8e6grASJeMS4+OISJukTAhNUglsiz2oLkc38
HE7kIy381Jkfr3F2fpbcdv1rSuT5DTPScIUj2jyo4IhYA2Af14UkTgcwRxwQOfA2zF0EWJc9KQo4
cF1hfX0AzAzwlWoyZ2exuacAqXFckPakOzbDwFfmd52NH7eqjVMkjl0L9UHvrvKEXTJIP1KYgQAR
ukTa/N2sRxoCdEu4+xd/5yebuUWcxp0CCD4Ds/xEaDr75Wh4TP/l/cyL5spF+lmnxPCYWT3ga/SY
TBeWNVTuSA7FRlR6N47ao92DghhwbN31zfiK/A23IfQK7tlepYRizAI36kGFrXAVR23IJGPliU/P
gKctp/fUhOwHlItWcvNm7t7BQcASeg4k9L314BP3cmmg/JFsDdpIIHJqggWKWJqDbRaZV/QfcBiL
H4Mdm0HEz9WutY7LKJWTYmK3WkMwzuX9K/RUi8cb47c8mWaAgpa32/ew8yEn7BfOGnaLvgs31hyP
fmJzzn8wEMFQuD9HgKT/BT6/JdtmdfBvdAq6RrbZiIl5xryTxEnV10RP2KL7hUbN0Kw9rkG7LL2C
kD44yzqPprGRHz5pPdTSQwTENIVVbgw9PlBeOxrBTkdF/RTMqSnSUBo5ZHDZIz2zWpXpjv6Cj41b
J+X99p9bZEp/fwo589MotiGlJx7R8Y4iJisRfBaM0bpZxfkb5YgIQigP1jDNwx7UmpJMzj97P5FJ
vCLV9SMbuN+rom+oYFCGzLcuHdkOHm+sfIOgGVaj6JATApbjnArC1IlbcA8U8ZapzCSmFRNnDg3O
IK+K0VFcfQDi/R06UvK+yyRETMWdR4EFh+yJGXNaLmm4tqSZVsUeOGTsbOpeM4Npi/68roELkuhi
ecC4+W6abGZnbennlMhesIJzUE5R4K3HMR3Dgx2TmvSR8ZeVm+vMikCEpLW/uC21wl7fxCG4Tsqr
LEuWspNP6XFEbYHUWkqP7m7PEwURBKwtNvDSPb5emH2ePJq/bYgm3/nyhYf3glmJgq+E7QzFLl/S
eR7TlrcfTnxrqlRhm16ip7SJtJyegCPP8wBhUOTDJlDPj8k948LxPRAWt/gd6D/xyNWf10G2VPWC
roeQpbAycAKGPgstaUtyWTziVBTAdGkAlBD0Z3pmK8QCSFP0grCAZ/m35JaHG3Ikx1ugmAl4kWfS
Wft9Tl84+XXNBKbNACx7KIVs7s61CplXvfp15hnVSyYYEN3gY1L5su57Dms58icJOfe01G74Wvvj
AgNv/pYwOo7D5lhkK0t24Rha9VtNRqB3R5vFGHdtdzU8Y97kk0UeKI7TtyeSzO9X7++SEwLocAAd
bQrZfM1HZdQyr7nLlwlrHGE9Uxa83eCiPdBwi1USj+TWyWTEqtnT/Jb8VuB/x97sekXkPkRfwOiP
zoRCS0VLE0kTtRl/qjDS/tKJATQGaxR6Z6nlpqBMtXfpIcFsn7c049M1DUQ/4lzdiP2jOafvFg97
x1e4NtDtV97cjCNb1p86InywumdgDaYA1mMSdLmZkvWH22L5kyfMCLt8p0F+n+1KYVXZ3+4hYBHv
/2602mngJVx5uDUjyV/ZFiIiQ6+cZTfQiJrXM+Y7fUE/HlONxBq06HPhcU8Xkatc0F1aM0kSrIJb
iIcMimXDbj1ddFu9DSDcXB7UEz7uL6+au4zBsC2C/+yHQ9qNPNszE1BtQv61RHNH+1c9XiZp9v6g
pIAbZ3H6rDmL6qSYMNe/b44CWxREbNlcn3+MYI3Gj+SZQwmDfTibA7WVw66DeFKG7u6PERKm3Do2
jBLzQJ9cH1Jc52lEG16E6h0Dn67fHOQNnKKxF7A3NBE0j7mFy88nhYzEnAoMnkDgVQM16YTryPX5
Kuggzpw1xxqmSBp2Z3xr7vvyCaBZBKLbQH62kAZF+uQfO5mec8AoHzD6EAJ9OciQsZUCzPNZFUqz
7dgVBRjrjLGKyEVXPENpA40WTMobI97CW/5I0h9cAY4XERScCJRH4sFvhFRV7jcrSvpC8UaSXpTQ
h2LX77MMVcIse6t907UJx1GEvzdThVL+ytOgD9bJHiG+D7YESY42NLG6mSZ3IeJkq3/vM61Nnlvn
F4g8hlaVoqLWYQjRtVJ1Y7GBq/PIxIETfAQyLEqG94o1PMiZE+fiSoPAtfylcwTZPMU1yDEnIMCz
M5eV0gKwnw3sed7hvkKAvMdDrwbIbCA7dQRf+ZoH0uM5sFi/FrZZ7J7YvREeZxSZRTYRrCEg8iz1
qRBgNWCMEb0EYbciJryJmgyTr+8BZotOGMunqQnGIkjju9ZV6lBTgpzLblK2huVC0Pr4BBHL3RtQ
iMl+58E5YiKDwnnQSFNfZvxabBrLM9ckh1FqDIIeq+/NmCjlqb/OwJxDLR/w9p5g0zQHMKne+aJp
Etd5lz66HsJFsj03AYOU+5tIiBvtU4f+sEanbT1zDbMsqempRT7kvrPVSOoZ91QIMNlngIWiFcfm
P3nXdc2GDRXooVPtDi/4/xDhtRiyv3wC+41FSecRL1bmi7Xqa1iPu5IfxIuwukIz6ICq/iyoXj8m
W7s/N55VTSX6nGLL7GAz5SGbSLUtTniFmJsaeypwiDd0PgtjHsHc380xhxbOCHrdPuz7mkFE4Umc
ZkyKPOhi426D0ih1VNlWdD29hlNlU9/zTxwp78/5dpP/VdsXIbSFkdmgh15Kp5VPYx7Ic8SduEZ2
GW7PgR75MnRDDLIklCpWxUPGf2mzky7MmogOq4buoOVwP4TnI1uTRvF3HlgpkdpZFCEwA9leYmGm
naTJviFXkZerZ9xElt9kre0utShzk9g9LLjvvTyA8IAmXk/guKkF3APqV3y2Bn+1mOgOEApkhBfJ
VOB7e3rxw53VBFIpXbwf/GcwRZ+ValaTQjvjKw5wrD8BRiMG5E9xcWl5gJ+gqEpZZymtFRo+ss4k
vwLuUdU4NS4FNmuddnH9bUC0gNUytchX5ea7li7evx8nP3jVITfMXpaKRTcgVemdqpzgu0oHHCWF
GXu7hBTqQrOCaY4Yabp6QPtcKmqAsYF4MFNU/nYX2LNfUYLaw463DMjxi9kxCLj+Q3O9WX8nkbGX
fHauXCGouvowsGBcC6EaFBVchOkjKph7ZeGm31Az/yrDpqXypWgf4YW7obVzwD+wqXRH1Rgnkg+n
qgs1ksVz+aKm0yiqlkM1NJXNEn2sKVzsXC0wYmaAuSohHP/gDcpf/vRB7bgN1WVCSSUAGn5faqh7
eoxbNZ5ikrDOGGS9pKHCHkoUNBghiNQYtjAHAFO7pWDHNv9Dz8zdPbfE0NTBqGoaLRet4TFdMKRS
YqwZDiwdNG5+Qhmd70EB3+sC2Ez89Hdfy0chr3DalKO6MPfGzYmy9ZX1NFSwSyUaDHUqUS+ZBVBM
H2PfT74GVEYRLSgfP7Gte5iLpIddIAx6ozBxltxatxliebMnrkZs8uO9N5QMzhRRKD5Ji9NiTnqa
9LJrLzBt62hprYqIj5ck9ZfZRrXVKlghY62Zv9boPb8GnXNPv5ybPMcMEJLK7Hm84lCC7FXuq3oE
zJIB7VDfHbtCe1p4oLBAzORgN8LI4YiZ+nf42d3XXNSu1lwNvk1Ms6THL9EWSS86wnK4Ue/mZCxu
4GMlRyt4vY9gEOd34YzwdIpuxN8GDNNqHGdLtkitZhiJoBZqWJH4PrHTN0yDlAaTCJHqxU/DtVjM
5du+fV9l3uQRZ0jGBqqXkmjiD9iyqkg4QQlJfasbtHxx2LhG0spu7CqXF7bnGZjx7zPAnFJUoejp
PHosu6nfpTv6wIRChZ0IXCbn6rD9WWzYW8tf3fzJQPNgyN7byCzjmNFp6hJc3omz9bmkoup4HhYE
27buQXmYFWKcS7g3NlRNhRe8AnHW0ZEB0oYLSgqUje6G40fFWnZ19iZgxcEJREqfOftt2fsxPK/M
QIN9Tq2ywa4/mIbol+YCz+2GGzSjRJ2IP6iNgjdTzhfCqd130wyJ+61eBqhlYRi7W2GUUo4onDiU
Wa/B/EHqZqlhAPDJ4TgfQT5byQJKpaN+iZMGlyoCwhNjDOEiy4NNRb5UiRgBWqS2LH19e4b/U5do
NsP8uWqBfFkZ4bVgN0xdTj5C9K+RSQrYLujPJpDjzM4C26YmkQsjUnjuATfT6eQTZWY865t8iBOU
c5oGAKK08ciKBWacihp6mZI6txzznQ0ZOVGrrDlCqNQrBl6qHTf2eNRdbmNxTziWFxPMDBsVyiQC
65KpaO/791vRV4PryBI5BczmkKkbxOQwiGP9MVkfZ/A9WvvWCNfz3WWyXdyXuXLs0ApMVNZkDaaj
EYdAmZbnq49y9ni8RWXZUi6j381xV//3qAqjTu24/CnHUODOxdTsXBirEBL8yChkRGHI85oVJuPP
PHwn0BZufl9Z6GwQqPpoUJt5BDDADneXvkTrGRpE+DeKkpUYnJC9JWzJyW1p+7O1p28ZeHeFqvyu
xKSeNB/wD8li6/lyK72SlHH5J6c3MKuUFQk9OKdDrn7g4ujsNJsmLG73zIDekaoRwbOAD4rkgyXr
+Da6U/WOKwViSPqUuxLLEnPb9sjH0ONa9PDv3b+556SjCuRM3yIgX6jia+4Y88SApH5ewCA2nQrV
7abkty/Rku82OcyG9w9+TGw2Z8cbaUcX5Cew6h/Ue+2UjRM2ga/FYho6godtIk/B6CUZh92oJHLc
7+2tRVtkR6AQhWxeevu4Os+yrOwrDgKLohQGfKBV1JFhk/78IppdMRqWwdn9Z5eN9VMBo/SRZ0jG
pbqs1ktglylBmm/b1778MoTdRyiamV14cYmCU71iCl31deZi2sIoqR7hEzSbjrhKQ5rDbUO/lmX3
IB5E5uoyVlh1Qt6GRTr6AmEILylf30DdeM/757Yzgj7gasBZvafZmLISt7r7CP5jeFOqD6gVruAN
u4zs7QIfCZVjtdH2saK92g/hQqSNypi/TCwKd4AR3OODMECKOTwRNS7GPUPAd29N4qHXVelFX/ml
MD+XWSUJrw9dEkluQyPoJhS7y+t/aeqnRrpuGEVTkgMaooqhBEe4+6c2QkA1xs7a6DsgmheMA5V+
C18z5SKyFQcNlATBY5SOYqk0Zv5LTZlzy5TDOcrON9U7o+CKu1nmUcTMAUrhz/pRYpkdv06SMscs
Tj30JVI0XnR/tw9mGwDM5mIFwOsTqA+MNVjjt5xk33SnFUhZVvupjenVGrPuizig2/1ud8jIMD2c
iR+IfxBfMxJpbkZ2JblfNoDO6duZ+xtYgEk7gbTDy60kkhsYYILTHkAKR432wHiQRFmlkORPWjdg
TuguKtUo3BMLHW8/1uAVWi/xn9uPGB7kxyfjMicLRz01TOeMEaka2klY9zJeZxgj4wpwjDZ53Vu5
Zkl++v9SFwWxnpPTDAizw+ks2MFbeBKof4pyG4jRJbd5aZpJcQ3fabYqttMYoCfR1fvWLBBPOmVP
uP+DLqp36s8YJXLCxZ5o615QU5KDT6w9pMMDW8yaMrs5ZwxgH9atSlKRS73yhLaGe/qd6x2RCazW
YdAgQB+FjIbgUBj5Ll3fYhQK0E9L/HzNGzZuVp9h0zwZoM9HBqA45n/VFsLRS0uJWhYPGGrqrg7/
1LfNCV03Nk+PpBSwCUo3SFMJLwrfeT2ySeyr/5K5JiLOlSB4zDb/a2++b+LgVFmttvHk1WkJRUdL
p4eeMBkltAgRuvdKsl7K+0pLuuMYr6sYT7MvAS28YRYMwCuFTI5cHPYWnR26wRv113/F01+035F6
ZXRBu94I2mNsZXI7sNcLPr2sCXkrM1RO4AoLCvyeZGVB5Pc7fGZCLkYnsFyUphU863HNU2Kku3r0
orgCaBrFw0hRpEiNBPHUZ7qW31c8cqv/kfHvwQHfnt2Kf5yW6b8KHJ2MwCvOy0VldxnJbxU9wgmO
+5PMn0eM50si4umKc8h3G8eowNbsXXsFg8IQX7L8Lhw9YLKxIFwVygDUdUGsqiGttnShlvx/19AP
GXJVJaD+sODCpiqjnJmB43yseY0zkTS2XtChlfaVBvSP8rj0zmrSEthXCJ3ex0qO6XWo2AkcLkWG
MF5cji9evrVfzXAOT6pIZ3DK5px29hiY728TAp0aX2voKvvEAoO4qguurl8AwhxiL+cuc+2b12ex
7iWIwKFTg46bTDx02NvzDXNa98/Y4JEBhQeuN04Hlb3cH59AtsXCO4VuLJ4QSpK389QSaqHAEWkB
vWNLE4mdIhn4ugszNy0IRfMS/eLhwiw5T4qtiuJ7U19JScnfSPtRRwDn95iZe9TdXnVwh7Nk7Uwy
ns4cvYD51tZIGUzZrClLDCJYZBwSdvdWd8z8Tnt0Z+S9DBSOsN246ole0NM7amZWk4juCDg03wlh
7eHOeZj0cdWdrr2jUAg/9ddTzOpF+NEHevhkjuq7THCsF4Sh5hdPzCu2fAg2tKf4Bbgr/cBPULyT
5XWZlBa9wIQodElalRagVrPDkkU88X0y/O05JYpeYwqRjsiqwj0nbNqrjlOfXeUNCmc+tgIRK6bW
ipH0G9TwQKh1WPXOciL0pnrZWBVbeALg08W6YhTZdumEUN4bf6d2T1cMZOwJ9lIXpAiuzdrylt7g
Q3hjhG7m0/LMcOH586nLwQhbm22e3ol0NmSy9SnCt3/11u5zieO8GJSjcHHhjO9V5jqWtQsho/M1
C0UgWPDvFPXkL1z+0zzCF74mai7GMTbhyc9ftsjG4NUJiLCo3/14LS7LfqBvITJ6SIriAnXVarNq
A1cABF6PBl9VkTYUnWSWd7FXAJuMjggjhEbs79kWlMoQz27h8rCf9YM7DjbuLWyMxte0xH0yGeYf
vGFEw3pKkBWioPT7KKNMLtoGG5WwoZGMyhuxzXg3u1ZkiHsQob9xAK/EPL6BV10lIAbs5GMdGcf6
IVcH/XR6ez3hhAc0Wd6N5tBs2iuFpo0FZYA+bU5KKhJZr8RauBMXE1w7fQ2m8lSkhPp67yrQ9utp
a89V5XfU5ASHA83Vf+NlnmJdkLEUjpULFwEyjDA1sIup81CJIhm3Nd2aH9Q+qlXjPZrsQzeX/UsT
XhWCUquwrlMvmY+riGrLd2ZzZvcppS8U7ebVoKuoz6MWXX6/vgQUFO7fjwzrtItuEj8crywY979f
vT5GvUqQ+f874RqYamrpEpV3h5sXg33mCx1Ww4jb0Ii9OEWzrayxxeAGQIxtBIvqleFmnk2rf2Fh
/3SIhttvj1ocCSqP/dHR0veNH36U1wBJRMNJn//olqLIaZKTy02scyhxgOXrOAmQ6LR5J4wbcSnT
wOL3jWd1bgB9PYhlLysA7ccvT21ySU4s5W0sMnHGWMaRsvEeMMMCsNo+E25RmwN+0hwPNI7yOUwj
CW8LP2o/9QHMrhHhnKsm0f1gUev2qlvS5iOMCBCyUrDG/zqsti5ydUoni/4eUac83QqTtcgium6F
jrxzejuxNNvCmJ9+uTjCMBm62Iptcoy53O5XHMTK1hWhgpLAcrPLzD03tmDt7yPvrEFvyvSIn8Kg
Y8uy1omQQ47MXTnPl+2/jTwS13o1aTNMjds116JV9BonGOnin6e3a5LcTTGuEJIhhkpN3znmZrg7
gebX3pLxiK+VnUQF/sSrKQZgpBwKXRMkk0ex4aypHT4CJPXW6ti8/exg8kplEnpb040/etZq2FpF
DpM65Pm9UNzopvbtu7tm/WWyunU3fr/SHkPxB+c6oBy6s42EdXbAuHNXyg5pNIE8KeQjT649ilUc
sRvrOV8mergPqr9wejd53TG64fGqeQIHjFwjPsUj87jjBiQpjsKMogWYxmcCGtNxpQvgwk4YbuyJ
NyOHHsoGyq0sVp4vyzYXt5U5INkOOPrFroA9eS7b+N0XC8tYEGezTi66nVmYTTxo+FPIf0z4O/L2
MrNQk41UBR8ffM60HvTgdttih6QPntBDDPkFOHkb8IhIHeQwfYQq958hDpMglp5vqB916BlgCUg0
ThWuvACDX4CktZjvLCkhep1HMdAAldiRmutxhB4s7wLAVYTuomlbrkB+A5K4ltxtt6ykCNRZGWuS
BcfTbjnjyHfnT8/LvMO3OUN+zZfLVbrkvAhDdYpUj4EBcV1pwfEHv75luSh7cvxJ9F3rwjI0Dnn7
vkhecrMojZxtb/NtPsMmGz5mIG25EDN9BHEDqEulrzl4LcVWe+I3snYOk5Nx7coaJ07pjCSFu0Ua
oevVK0WfaWCgkYj242QwRiBkmyKrbhIakE6wkytz1+GcCwyNhlwyRNJnQXrXKAmQadIR4tVmoxao
a9cGQAc/oEVme72quwWKnY+5cYKmbKEzoc2Gajo31iE0YuWwlQGXdvPr2UgRTmo0MKdKhYAxqXLM
J5PmIa32cckYYFMEDx2KskrTQBooIgHOYRb2UN6g4TiVEqPMh4IEOmmRcRzvugXsBmOGULiYhgHr
WBoXQVbq/ZNpuMJ1e85XJSY+GMxOk0w+GM/xZ8q9hAlxhobDfcqNT4q667wZHgRGjTdV7wQPbhRf
kJA8dgaZv8V9jpA7WWg8y+99cxj/X56JGbof7fuRUU+wdKsEVYXj2rhXI+R39btnWox9/AswTuLy
6aExlpKIEzPQ9gdP7I85VbUk8QbF0Jk9XfCd3F+5lp+PrSvk0YErluLeke/TA/8UUMensHh7mw51
C5jwfd1oKNLPGPBxgaqDC0D6N2RXJEQBK2eCRB2ZPSS/vWUnWxlRymySLk9bIA6kqk+ScWJmH+BK
9Udqqll9ugfpJ+IZr6zuRuSmb850vy1t45HTpX6Cta/nT8Nf9wW1wdlLgsbWM79dSQ31WAX6Budy
qdEaZGv3AWW11smX896nFS8+F7W+t4PsDsgEE9Fb7OyaHeI6w1dS4xrMvEPH9pQzBi4WiZpLVXJv
rqsWjYstqhevEGS1H3gUQ/4cZ/A61ZmKF6k9eANHEuNrGsHOzngKqt1H0VeJFus7iKwiC3UKsWmy
OaxmhmhaPjTSm7s7ofNihIeAnAO2CYs3htHBzmlP2WB4ACGl4rwQ/xqN8gKNglP38MiRtV1+/5Gf
Odwwflr9RcDIiaEDf8ObRc2ZWt0SgKAmUzV1HUwXDqY43ypMApvYwjkMLKVonLJdy04YFEKASuar
cSwG6Oi9r1mx+usQhMnr18/sIb59icz+pBln6ONvWfPBB/IlF7SNdEGrDFO3ghS2P7Fc+LR3Z3KR
cyT/yxkkfgLTD+vQ7InFjkydnGbL1dNMXvs0JNyRWI1cXd37y3eSHb/Fl7xKY6s2+8rp7Pmd+5TO
7qxc/Uh/FxWA7dvYF9aOnu7oxxSEU5m/lAhInvkCStKfm+fxyLvI9JsCOzozwKZ73iNKJhgZNxOz
U+f1sK0pkiJW7+q6dd8oHuBS+dlEQ0TdP6+5M31eBGRe5c37a8y3VsIG6JvZ2AyIqj06xZhGbyIw
ARxrcU2mA2Gc2dYdgQAz+kvC4eGrqFIVR9DIYOMPz2OUw18LNvjwY6ybM8z0FJTXIatxblNypC7x
SEn1Lht3U9GPZ5wdVKpadIMRCOnaLqnza/bHPHYfvgeB8EGp25zNjHOhIorNvc5M0bk5gF588Mwb
TkrKlahwcdQcoKhbgwxMPwRxB1sl8nbTE1d+c7gSpL7pZLlRDPfl/4GLqL3xAw2/OCH5TKNGcaj5
BnBPaLh5u9JrUOoMWL35B5IKu6Eu6va5hXZijycLKP0g4KclT6awJeQHUFexbOz3jaiNXTHIJUCA
vSX5iYU94wYmmLwHENFGDMSqZ30c2Jw12InDwOgoSReKQ/IYowO3RgdNYj3fxw2zlMy2Occ/6t2I
1285bsuqWkwLseTIXWLQ1JMC6FiOGz/aJmTcHKWfDYkW8sH385FdQn5z6cfueRyn/S8C5I+1bF9F
37uNCCWl5i2Rdq5fJ0YWx6ieM0jErJ5m1VG5DtWrwHgmsgpoCPiyQH41uRIKHvKA9s/nAAS6xtA5
Ylb3cx6FX4NJ4ZGa4BWk/ZjF0FqoT6ge3FBshKFjBQPJVPhvM4GJcqLDb3dGBgywiXb5IogBW55y
OddSM/J/lDw2ZLAl9HGk7ZS3oxOzk1g65FbeuyDQu0YuijSDi7JHBGxYT2Pv6vmOf2r9z6OkQpuE
qCd95H5Yb0eUZQRdDx6pvIgLgG/5o9/QT8XDVHUHNfcMkLxWJaMAwydCF6yK/EfXXVfDMtz6WRXJ
0pcr3lind4VCi/264l51Mhew0YIS7qgKgXZEuHpRbvANwNztvBg8TEdM+OxZFOGNJNQOxB4aE7Yf
nSZzZDdhBeUow5swrEjDjg/PB6Swev7DdRH7yjhI3Gnkb8BUBO5Pui60cpOO6MnEGnAiwQeeVuqT
1KA/+C5UPcgJnkB2h19TA1aigCCFsWn/tbGmBfP3Nn1J1VKJhjKtyN8ke6M5sVRLj3gShfP5JY/3
oYKFe5rrbn/Jra84bt2qm70l9+rPzKj+R9/EovidfCXcZQUqfNtPRJHe3AGgRpLeh15Au/DcXV3B
NRPojWTDdHYe7dgn5RWVPGfCinphNyH9OX86z22RQlOc545wq1+fzwlYLfMv5PjyhWjH5pCZMlPQ
Y8Mk2hTnK4V9TO1qbjxvlQrgReUII3QX0+H9sjN//4dikKQhaFBnbh/It+wG6LyQlRn9wUimq15i
Mv1L+u4hjxLJYIIs6lIecPijgmkNpMO+xieHo6a09wGIM0E1/3xAEp6w33hLJnxf04VqUyu5mkod
zQZJfPr4+bFvGt1UaD847f6YDNf27nYwX/BzCUv7LmW4o2Bdh7NVDfjQuFkT/uaQGtszNhxRraZ/
5Dhf2SletXJNZJ/I32I4Cu4JNGFlr5vvtJuGdv5mTtnSth1zp/7KsbFB7hYIVkLswSMPLpMyanv8
Tb4S/0f2tkH+2wQbUP0RV5ftS9zm3J2xy6Em/skZR0GExonHhKeTbiE1GahpOiywS4KbxUCtoNbu
RX+nc+wUqK6aJw77zWbIdifI0Vr1iY947vY5uF02p/BxZCcq9fRTvF5R3jEoAALyhK6KYmt7xag9
5zBoimvIcKxO00Z/EsDoDpamM9bygt9yRDbKZKmMVPBslBxLtl88o+i3IYknhuAmOpM08rvP6sl2
oRq+LkcJjhqoXacod2cHnbl3xaLnF6T4SnLIgsxeoTjjhYy/udDVI8zSuskp/C6SM/GXwvGrfbn3
ol8JEcxki7xCK4pkUp/rlqGL+tCEQcIrsEDkAY+hkCGPWV60lZmxvsyivBTpQBuXnsGfYlNE7vzX
bkFVE4zPR0hHVC6nfTl3II6PxbBf3WaE/TBrXImPzfUDP5SSx58ams6wEfsGoeK/1bPayLy8pbE6
mkES14M4fa93hRtyfNxaceq/TmH6ASXstlY6tvH5XcctF/zhmNvqEwWnpN7/PVBeHGLn+jgyTn0I
mhG/ybGMyH+sMdQbcTAEZgEzU/WTE8BOddtAtDNu+ntWbTIEKUp7Y/sDDA/UyEJC3LucV51buNaL
KhhJ9iLMGbEBGF9MzecuJLiRfiZJ/V/u5k2K3cTyGxcmgfhJtMvVj5Yo0AsZWP3eigTTiI73KgCX
o6YsY4AUwI/1XJw+agbg8R+By1Kcx1WsZkOSPDDQPd0v52ps/KB9CguP72zogDYGRQQULc7e5odU
Gr+8s51ArSwb77dnPuo1CtKTzeRurqI6kon407ae+Q3M4AR4gwa4RPcPih1MIlf/fzei9a3BuMT7
DZxpCXZjOsG727c9HsAimV9ynHqjKIsr7SDHXhjvm1YiU9MjpDMepibUjo3+D/fZd5VpdF98Inon
PJGTkQKtJpDCNGwyyR+7aS6XHILWSJzd0xEj5IvCLy83y9AglgW8knyFdmGS1T5G9S3Gbuu4G26Y
/Oy6nEGAwEh+7qiRBtOuKM+R1g9o45tsAg8O++LYEljXCHKTI4GQ4KnMCCFTHCCqkmL6XnSH3BoL
WLhF2o1Loxt7ZuDtO2zkS+srddWk679bXPeHhCLmhupRFm+09yXng3wHHJaTN0caf5N9seZsMIg3
pxPWFnPmMNRH/scByuWdf5CnX6xYrxzcmFyv22lTOH9DYjxVYESRG2IG7DVxHRBnBkumwFi/cqdJ
FtWroJZCnDH/5IrYjbqr0beq79R2JBBzzs/Q6sdjrdHE9w73/izT/eCETW7xzUmpdUBuQ5PZBnac
FcbpbhnWlEfXnovnWJol0an9l0/r6olUEN+ONZ55q4lSE52TFXZzyse+bUi0wvXdvVc+VEL6ZQQ/
lapAYFCfGngbZ2x1YKff6AOUjLQScKhD2WlQLooi1/A/EGfjsYKzt96mxBo1nUSW+X730EDVXbjC
oLVSJTu7zvox84WxMbn7v/b4qmS/BZLvUfwPO4Wd8jc19KJu5Smq4uagDPgWbUIWpQomzfDzWJP8
eGcIddtOeo16z8qA3KdEDkk8TLfnpgT6yFyYwWp0kDaBUJy+/qZvCTm0tpToEl1hdcgp1ABe899S
s9cF0r6lfGGGDnls0X5PLEShrhQbwcSRb2b3vjtn55o0A3C4y8GMBE7wVqCivZ/Kptvz0Dywi0yc
GFNu7D6jQ4zePQSHznMNgX3qBxZMZMh7uQ0JKxjJ2l2s+j1cilxBvotgefckdn9/JpX+SXnBulYl
DeouvwK7FCimcwAJonn3NNb+SVRN1p6PBrzi9UEkwV/Mh6Z7K75LcRPIgYJCDmuCO06/kBAJK/Xd
ovaO2dcpiB2sBVuxMKX97kTzey/2JjwdKCMjDZTMjpCt/1h1aeKIxm8QQEnzLCCZtuiMtJ7P5h0U
2+mPLAe/qTfoFUYtnru2bYIYzLFKT4yxAWBt0Ca5g848/hapOPsUvWaxBzwW1i01Yak+VdG8GX7v
dcb0qEzTgnGXAYxZta/MOFJ+IgrFz4aLDYm7sUlkcJUsBRlVMJpB/f5XhoY6A2Kbl+x1roRsSjRQ
EvueQ7lRy3daUTRgpyl9p9siThKOEE/PsTV7AzPf/DEg2vN/ZwYmqYegaxBo1A8VevIdl+gp/Rsp
wgFC1hf9aDTr4RtYsm8ZHMrYTOiaP4nZZY/dNa2W1aj/KVASYhqG8lyf87brZpWrUvF+JEslIN4Q
RfUF237Bu6jL5+1AMJdxcTeEYND8Y6lWJ9SJnfM0E6wjRk8p1ZQMsaqrOcDIOWBkoE9YxTjM61+y
mHhN7W534HfzKntT1xVk4QVJ0sNUezvMLOghcCM+amozxmexsX+PpnNbzBHqfGTa5IpHmnUDg9Wl
p9VPaB08uD9lwe2yQmo7/NGKVAZoEMBUYKD9ciqriNsy6Z8byYernYhThQEnPPDWa0B2d/NzczgM
9JoZ2ZYYBm9ihMfQ/8D36iFA1j44pD/H+dhD8lctAmJ83oN2INfiNegcaO1rZyyCDifxFJKouVKi
0ps7zVnDQzw74i+etGb0gKrg0/yNsHQanQY1gPWgCh+uVFIb5snEE4bRJioQlFeI3BfiZStmAtUg
6QDQvKqU9MrrBUsNBhhqVqpBZ2mHFodaxIo5/Qg1pkNPZb9sz9oykugSXK0XSrBX15T6W1RcRTS5
e+xjtX2FB8ssyv3MYO0SbWkVdstjntTrOTZ6AhqqpqE1VnLovL82xuktNumRXS44EiprSZb/MdNs
zK2uCjkJyQ5Z/F/yfDWOyPXxkyp8pAn3f12QhxfXNu9LSI1uRpsX9+DUUx3tuU4/axCp3rQvfUX9
RnfvlfAfFAA+GM+YBXm+SjpZeBknuc6vmmp5kyUWzMsPJGqjGO3IAcwkmPh07MHmrLXK0961AGx2
TEcvzLms6PekPVTbY6gyX8w5g9ioyOGtUrwz24NeSmlAfy4hZVnLUFQTsHLJtE/7AJXzXStAYwhJ
9SyvuYmpPE3NvUbk/d7ZSIOu9mkD63UTAwv89e6Le+KPhgXNZza78VzRE8aHmhNwenVGvK4na+WN
eLoLVr+aHvEyIXYcy2tlBMqNkC/r/pwesfHCJI6W3ympZYz7JUJUrwnelb0HyKdJiOmJyru/I/DF
Y74PhlBpld8fnWt55wcJqLDcIeZHiyithmQLgmzVPW5xq8qHeA/wTQVvJ/ubSo2ek5bSak+dMhVY
0b8kMhumuVjtXGNKr91BSyxzIs7S++gltiVH1LGHOqJOWX4OAMx50d9tdEo5J2S11sGNeodpdYPx
vnConY/O/bPSmKnDxed2yK1nooTeKBrNwuloX+U4HGDYOEGPsYc+bSv+KdUCCmAvWbQJf9eLfnzG
gF7eXGKDaHLfc8A/ZvXwf3IV6RuIWIOfgS8Nkjp5Hvg3d6lYeu4CNQm2Bi3UTbNHM4bMk4QB0sbF
cfqT6s4f/GflWrGPMjH92WZf0hCB9o64xHGGeO/4DuOPk/fX4HKwKxOncmAgS//mRk0Ml86qekpA
vzKyPol0DmwUUEBLFQkMN0rRv7RKcIHH6hd/XdFaleo4vlsxUaiYj9qJbEtboMg1NR+a6lD4gSlq
A5Bgy9rr+UP7/whOqjK9roHetKgwGS4/tgCEn99pZm3kM439HEqasj+UksmH2fc+Arsn/tpBRzis
AHCbSwQwDJiiVKOlG5GsDlckq6BSLKl+h0YzrpdjjwYpz/YwAN9R0ZbgDK1CJ/ucrYJaBBsreiJd
Dl/ETbZpKRXJFgg2FpnjdY5hDy4I3Q5apNciwjcWvE0zksjxyFeqvdXWuv6jhBYsR/QcgINkSfqR
ahSjOVZXshldBv1km1LCt2f/kKpV/bqZmzbgdyY3+Yix4ochYJmNhSCBvrRqtxge4ywoGfYncyd6
99Sx2WZKQagVO3Yw9zqEwJLZyDhBHUCw5gJsIVe3BIwGtO6sbku0vxFgDCkrI1DZOWTTXAU87jzw
cEJBdy4TCRo8JGefIHRHGJh7aVjdQZp2A0EGr5jA2ZL4NCOtUIVtXN/W29H1qIDAOzjhf/RBzL2o
X/pUAY9ITjm8Bz6l9W4jc1QLYTOHniqb8Yx5T5j6cqDVOQDlrW9a/yPEHiAkcD3TaQYGsTXrRE9p
cCDqqVUr2+Y7VF2/LTDmiRXuZVHjUfrpY4KWvam7FzZdrLgKeeQB8HW89TTHuCQNUGz+xxjvMiPI
KXQ1XLyi9duNUCfCdSkvhYANT99j3y1Tj3TGjBVgyEeHGyCKZBxk2FRtk7kL9YFLQLJBgi7QlgpO
Kn2LlckxiAWeLkCaJGab+wUkfnthPEfyMK+b68m87CLiwMcXLy5Bc5OmzS/IzBqFCrwqAkbsFbnk
CETaFlw4INKUGY4k1YUotmsYGmEd+OkWuVjyyzJg1nU3zHkD0AJ8ff6YxmGqnGlQH4vpOT+Am5Iv
YEUTPuyj7TcQY2uQO6Db1apqFwsg8isOq7EJXD7RvwpAd3XdLrkNGsRESKbpVPXtko3gfp9Jj0ue
+wy8XRAKBs/pDJKTB1zNwi4KErRs0Ed0QY4uJR+rC0v2MoVS7VcL1j2jnyzZ2pNtwvUOzSXlan2r
+Yt/DsyEM+3G6SkseeX8y0HOFZUdZ8SS+yh9huhvmQyk+5FzlyqU7w3m+7OrtJ09ReHIK+GWUjPp
1IY++he5hLuYFa6rp6sw/5NAEwLUAghRjKDwpF4Z5SWPMGRpki4FwxRQcroBmNBJ1HNd39FD7P14
/vmsrwg28NjQf0NUyz8rAMmg5ykO503TUcHZ87SkaIMR5s9PBrYqADizOl8sl1LKnmtfDv4ZLasa
LzwrZqk88SXt0i9ygEll7kquzYOF2eZ5+3wB5G0BNXm3udystsP3pC1TVAZVDUSGKRiSKAb2Ll2d
c25RkgKautkAIfs6HflDJgFAf91vawck0tNXJorkQPCGGuey95q9GycFQIml4ETRPSpBqQNWIS7Z
uSqkw7lk/ude5qHc8N5i+QOaOHN+AKm+TTFBoJmYFMvjGVFKfGYCeW3zWWiYlVPdI3QUXnLW2LFZ
Cf+NcACeEIh81Hs3JdR4VyTURm1Qa05x36fHLPuOcK3V+QsF+T5ZQEctGiKiG81PAml6so008uwV
oFGObDz/YHqqX9uJg298ZIZo5Kh87VfQpqV/Oy4xKc/cOTeBHDm6RHbmgOFlrOJz8XHSIeiBpuXx
5AH9/DbVPdf4WxGSVadVa6qxfbkccc1HGOP1x+NFFEZMmY0nSe5DdUJcs7GGsA9pLANksGy2IQ+S
LZdpyOAVb6dC/iEGebiSAfoadC0Rbss4ZUDvaI0A4rE6htO2XGKJjcWlPelUhBNERDWRS+00FBQ7
z4GCDWy6UaDpUavPx3sALry5qsJ+NEEQl/1v1NaN09g6muqOiuY2dvFXQvxtJoHta+CGrPpYWNTB
mGA1ZtQLCKuXdAO43S4qlCCWWnFjvTBQkWo1H8vRQltDD2eicF6JaGT9R1rWHoOPcAevUFoRcvfa
DdgzfOWWCrZV6svN2SyV7/feE2BGnUPZwDJi7qtvSEE2DhNFXgkFAeUv5qBojk7CzHWEOSewuMQO
vglvBbbv6oGhCLrqbqR8btsmEroOM6jG53Y+degsEYrTJdBKYQUN33jWt5QDbwsINTWeSqH5PEEq
ZUj3GzlPwUBOikZMDdp0l84qYdStkC5ewuUo9IvNlLDLCnsee8RUY295uLGW0TN8lG4BKspUuIEQ
F4hnFrjy8Aj8JqgychpEv08leijzzykaMDnVq05wmNUWObdv3e7PgTIdm1eAoj5yKkhgOul/tRNW
EvzZuJW02comHPfB+8yf1HPpkMYdzzeOcUI0oLMPMWgHKzdtI6kCbKBUPeZAG92pLwYUvyfJfX42
ZQu6uOZWmEu9grcPDXOJVikfvftuFgoh+G1LUs07NDpvFuxO9alEKOhzG2vXpZBdBxFvvo8jNvBB
l1dzNdFGHb1DTLYkCvKOgzlasLH+Gj7oPVJaKYANbK+U3dZtw36SMa0UwNqbLi0VlG06Gvcb63vR
tMzFzYdfj3n7V6vdbnXwChPb039JeW3QAO8uFLNB0HsMU0G0aXCEVsuZsmmaJy3eyTsNz7oXvrZ5
zvjk60PZ/oCFCLg1cdX/enL+rjpo5PlFoTels2tPpCaOvf7bQmB4cuoLvf/DOK6H3yy3Xm/S0OLC
dfIQ7VxHWVk5R0exrFWt4YTk2n566Rx36hZeOMwSA2dRosbFVSL6dWpFCZeXVeatwQVPJxf0bkHf
e0kD5ITGsvLq3DST2pYGEHIeV6DxRKxkoVG8ROIrY+DWuNqqyaza2ZySIjOBau7u2X5WR1aEcyJh
2y+DY9AdLcX5vHbcAJPAjOzyp1fFbOB6IRJa7HnG3RMQvo6/nMPAlxz+/O+dmyy8dfYc6jctceHE
jfK5Mkek4MpWTUWgivD6rdSOT1ygpQt6IOWHksO071WfWEJxV6WGwgCBYrpIm29NqwJdfs+S1me/
oq7kk22+y3ycB5zW35iv6s0ee1fQEVCktdpg35a+UvNExOTJnpkMD7qqvLNO1Ipr3WGwSd/BqMNx
DW/mHLlkMW6AUHhNjk3v3IuWMrXZUX6JqhDxpt7/t93PLvATOVLwOPc9H7+0xhN08gSN3gez3onm
WAThXjBJnYID40j00QBgIit6HnmC30BmAvFM45nrQHfVCFDfjYHxyRhs3JnYUNn5KM/SNnSppMuE
nmExPAawRx3/Mg51N2yR8UKGjtkr8e8L0u/HzXUd37cUHdL9d2tjRwGkuZ03fUMv/FscXD1iOTeF
rplMOpuCYZCymrZIA9eNQ597Hqe5zsCwkuuaZHqMARMhqkCy9dK0691A/iJ6/aWeuPUUc7jBrTs+
1hxi8q4/Pbo5wXLuAHcZNIQNFtFJMbUkPoVXI1r4tGzqK3ZXTRflI/bMj6jrChM5sGZ5uRUPXMaW
AFbfsmy70tj8ZEwG8c0husDew1TVCOJ55BhbMs2/kTYXwIvZq/yDjHbnXxRAyVXf2uqhwJpTdiTE
WkyBSLgaVXvUtkuMt9Pbv/MqQ3HCnTDKO1MonV365KUtf7L9cYPdA5PeL0b/arT7x+MoA/S5MQpd
qV/UuIAytkdFNKPnXjGOucx5wogFgHKzzaBcG4VKyB3e0F/WzVTlB7DKGmVgJAEStELy8VhjdoYA
X87p0aYkVOrICpOBEpzuMEemx/syiE5P+iGpA3FdnEYAFsjgmBONWfcuPet53Cl+0EvyI7PB4Cn+
beUVaD7szul5IfVSX8nFbdoF5jCZEdIkdYUuUyu1T0/ISTdMMq/lujvzlKQymHjQRy1dBnFJn/r9
MVC7Du4QevqeImWMCznIpwR5v03fcJWJzaHjChvms4y3yD6IqgD3Av/YjEK/EBFvR9JmgM6wLLGa
lSh1pZV0MHpMx3Jn8Q0O+J0676TGGe7qaxtcJPyH47TmFsNA8LFoTxJWUmtIkK42xJMvMniok117
HUecIZ3Lr7fzJtBIaMvaIlWechkYyAqsd91u31zIV05giheXcyAbZQp9L205m6f3HqNd/lS959Py
rvzwD7NCAV5RbKIOtMaZGyghQJFGitHzPDsaIZY/zqJUm9wG3F9EAwm0zokmP+6lT3envJTC+oi8
MOMjg4jvan3Lk09rBNtwES906wEaq4Yo5097WbVqWIUIIv3Sczt/Rxc/F+3+KWixhtYeJXre8NjR
roEQ+AkRMbyIWAs/RaOg8eUDfCyGA1LoVxZdfVXEyhWInCxNc5NN8+mR3Q48G2CfhBzsgx3rLdT3
utV5OPwI8Oo0wu8SXz43KdzsLDO5ev/++nOL2BxGFdH0EQBdi+2w0a5oW+YTjFhxGEBJ54f1xop9
kclFGUT2x0w5EO+UJSdnkm4p1aWCP8vtZ7aS9ABOcA+D/R1h4r12IfSj4Y09DFHwY/pKxSIIl4QU
lC5IG79/lHPRHW5kBc4kOhx9SX0z8OkhUAWQg26M5TNuit30M2fdDyIN0Cnawx49OlSLVLhmTBzL
nhuDDsKwYr9IjLQElpNZJv+IGYV1qJ31RIXrN12gx35VC4GuL5IEWoEBgHHl6OinQ/mq+GbGHLoI
EVFI/CT9VelWXuAA34y9UEZE/vBDOD1Us1o1Gb75ttnZN50HgdmGp8zaQG4Rcf4xU8nYZZfzJ45w
NTXHpNZYxEf05/ksmuKL6tEGDdUdlaJF1aV13bWsqvFhrkCQRUfYISSSWjsLgsBslBpcRYOQ9BMH
ZjjNlFI9fMnzAmseRd2HPxfWa0dhhiR1p2pIanWnxHpFXX8U9zy5njZ0RgaFHkICEsk9qAkGfL72
WkNnHGIX8e85aWdW+5CJxJXOy84AUytPLMu3/XeyxjC33juy8yFX/F45Je5rd+Gb5bxl+oeFghfl
/WBlsiu06ekzHXDjVcYfH/9WaeCqZsrY8YUOrC8jKzmc9gs6D0dCnBy+AYY9MD5itBY08RZGNC4O
79I52Ca0Un4o3OrrgSVaB83uSsPWkCjH4E/W1wtP2VHdZzQFZL4Ss4UehVv3Fuy+JsL7Z3Rh5PJv
rkAE6akmrVCfkH80YYzat2y5d9bCct8mvHKsqIda/J3x8j6Ikfuto6G8Aeiz44kOO4Q57FGlVtXT
IRjeYxUTZ1NGoD4Nbbxx/jtGiegsJAWN6ywKzyXuDfTtvcLskSd4ZpH8pcgtBuZjyX1AuUwntZKW
DP6OCwlMSUQ77gJ7JM0G1CCG4RSkVqNpn0r0FCwLV9se79IHqiNpUP5+H+MdLsH/lzu9N9uFSuqH
gIVgEKqTx37COQh+YmxoleMt7ootMQb2yrdbrxI8TBXDWMI1fTMHAR0NTf2i3kFg8oxRwQR+tOGg
h5w7z6o/ScGYBUEMGzl2KpSfTsKJqTxqpWihbxCTrBXFKBHlgd2dq/L3dr7d5NprGVP9HEZkGQRQ
KWuXhetTbtcIpD8ofqgis6UacWg756AhWpHTb1Y/ew/ygOgnI51Dqepc+dgd0aghFrGD2fL7bfL7
B4ez7TdVXyAdzgQcdsSHNhyqLzqdneCuL+Rm7Tecjgv76vGH+xQ8Tmv1h/k4ZMoB3Rq3BFSidLHR
iD447WvEjqzrAIqsUWFtMYmo9WF1WxwC3BPh2/Anpk9DgKO66uDCjmaN/HFpFrvzL/F5J1gzyARJ
/tiw4E60OE4e0n9IsqNMfaCI6+IunpNtt0OkRDmt0qHZwaXpaZZ05hMI0PuZmQ8OaGNoruRIAiMg
eAqzCwBnUc/cef1xwlvDAKJPsz5MsDcSEIaRXfH5qVdmyEZghUksAw8twHLSLQU9ADHJ7xIaZtxv
3naVICi4MLNhmGHXSzqUow98OrWiSXw36cOFhCuqzZ8GuEfVCFoKhMO5pjweIcb7PuLvbuowc+VW
dOgO5ALZ2tjBe1xLeYCyqSqGyAQME4eQztUCXioU1jCKj/TdEK8hqAESo6mehxXp3sBvBjzvUgKQ
s9AuUo964fB807nc4UmaczOYMQphjv9dBKzw1bJRJme2Rhgu7yyWThCpLENbsIVgGw/hpLGcKqB9
Ap8yWPonK8IZi+PbwQeLExMlGu80K/M1OoAVFIb7U2KT2UxN5TIyIUJrwR/Mgz9gmpO4AaGzLFje
KIT7vZttScqDnEVrdfrgl0DuPW+BQiphQWBLFb0o61VVBKyuKRYYLB/kU2of/A+qitcfl1xMd8SH
LkRwq9OHowdEUpDT0Mz7g/UgnW7BFRZHRKzWtpXVvbTWDso1EKP2IBzUsavBdITY3sz+a8vOlX6g
l7YPCzZU67dBXitre5lSGEW5OOm0qb+HzEGw33c4AvrLG8TqO3AZ4wL59h/p4KgfxrEEEAfcItCI
vRIJ1iDv5EHX4rh2qCW+riJXa2miVftB/505+WnpY/YvsTYas2XKI+nKgh5c9kCHIFKQzGOnk24F
7I5io/CrfXV4AOkB/hukRcTMutMS/rax9ErfosJEAgH51OR1xbYaUeIc/OtjwSF55xWoALedoWSY
a60YQYuUqwSu37192T1mrdQpMNJruVcw/uBiYmvFyk0uJII8NfShplOFquY6LzYFq8DqzUB4aUC+
+IjBPPU80MIRZt4MuO0wemsyrDJFuAVxQbN/0dO/cI1kbxGkfJazetLYxxedysZllHTXCSCYBnVX
b8A6vX7LDMA0ux4IM6wzDDe8PcnuPoFQ8cvhUHjMy735wnMwJ/0/WTv9jtz8Cp2V704CaWbVo/u+
IRwrdAdHKaTHIsjvXNW2Zx5+xxFfotoM6o4YWzmoC0LicDI5KtaCaWO9HqjnIqtVGmN3ZeUjklBR
Jimg+lvIW8VhNDNJf/Qu9CzVuZ6i6INNiDon5fYn/d3mu3Ot5XFi07hgpyR3ZCukoysdKkkM7OuM
/BfXbSpHCIitSWbkzl+150dOHufR7igdPFhUdSdPbWl9NXRoxj0wY9IiW8yC738v02/Ccg2hN5Xa
wW8RNja2NqWveyrvLi1vNxMuNzC+xjYXvmqmYdQsmegJ2KtRGXTlR+STlAvVMkBRDsMexvBxmw/H
/+lyp+eZoP9cReDWzILET2AWYuZ/5LSHTrJBYGnl87luzrn8FNE4Rp60r8eSgZL36FTuqy8vH6xx
2FOgwMpsShGvApPiWvKD3P6y2Po6TwVHQZZAQtlSObWwH9OMVyj8tlQkY3fKjXa42LGfQc82uf7m
MeRnsPzgru4tIiCGbOXkdLj551ExPkS8y6QrX6e6Zl+fkpcgOxsgr5GjjU3/yZT88i3ly5G6Wmnf
kfHWXxGrts4lf5uf0J4iLcjTF+peJh+kW5TQOW+DqsvWTlPy+uJ5kHIirlp5jDQf9VQinUz3LszL
31f7SxPgkURFgYlR1MMzCQJrVvurLeLFCClwcHtQgyVypwf5chKXwGO6ioS/5wDdwKlYvyJDMpn7
yIRLQIk6giwgMk0uugQVLlbxKgsASNr1ktLZh9ld8FNWciub+OtRo/s9y1OhjbozJhMHxCqC30S5
pga/8UlUk6TNy6tzrpKXbCueae7LXO/jqKXJR5aq4rsWiMkbt/QG1fwE+RGiGo8claJN8Bm6mC1t
jHN+VhWRWiqMfl+hiNUoyKvc241PvlrOibpoq20O4vQu4qSors3I2L5t00xfdSvB4I4RetgMSeCN
WRapYee3nVmVAQwmBuXhA/TeG6rDIo2RbE0lkWkDMQb5S8N0zblk3W2m5UrCvGgS016Wi0JONlxg
5Eft/UDh9lptKejQFnJ6oyBUn3X8f7FXi9VH/WdVhzbYo6JaD+Ygk9jjAzofzHUu/64L0ZJi+drN
Z8vOii4lbdREwHbm38GR7BFqvTiNA94Xba3L5v072eE6QPCAJrDgD9e9LA7dFSkOiiENDyXzeyCI
cQmeEB+uk3WKlEqcuXTdrREtD5r+HKg7rS7YDpZsIjetdx0eKuBLqJ928HdPzkR0egrKUmEw4fMO
QzQ2nKOUFbgHryytOnQv8lK0r5PANt9zhv4dcyePGiAifUkHwE3FhggDAQEhOMJ+3EDix8q5Aod1
af9Q/K+zr8YOOQ5TMRnhhk7rUNP2jIF9I4H0FtCbqgKcb9H+LxAeAg4LMiJhccYxMEVDaP8X5325
0PyMv1S9yX1+ujc4Yp/Iu1bd+OVXd4WlmqGWFzz9JjZ1IDhlyZoWwdo9sSGoYZm+B28v1fkVLwkM
lY2ZPj1dCc6TXmgA9Bw1UiZxd2DDg418kWDJCpoL3vasZ842RyuKQTP2GuXNwUWjVp04SuHRB5KC
7gUUjQU1dhMAyjRo15/Wvi8QnH/FPBqn2KpB7rzV27ecCx0NmyXPguRm/IEYObb8RyWoo050HWok
p3Dqe9BJlM3etSirBA341yCfAGDkf9d5OrXqu2gW6WrLWp8EnAHYvfR6AC7NSI3KIa56PhtRCC5s
2ncikEwIrkcG0Q+uEkor7tOil1q4+Z9rL25UaOj4hv82qutMRmANDt+8KqwKCV2SjCnYr4JZP0He
aKsjE26JmOj2eqC/Dft7LwgtwHIPuaWKmxc/T8eaX5Aiyt2Wvoy89tyUwIqTPo7aGP1wuPyN79F+
KxKqWrb6NPQLhJpPgRV47p2jEpcuDgIQW1IHBtyalv9F6rmQyWWOEFQCIQyMNkS/ZaHnXx9I+tlo
WxkOV4vou9UO8qFO2blFImA7gvLxhVY40NRhSw+1eq1rauD7dXzddNeCzlncK2TMpu+28pTWyJpn
1S+wxmujWLVlgRik5v9ivfrvqXJBy9PsQ+Io3VlFFlhBkfwwAiX79Gtx1wL7O6vUql0pqkB1AbBX
O4vM7QMxXiKQhh749fWaX+U6QMe1hTFK9AOQA+dWAeQcT9ZnDbf3dV1uhFjXErGYeeY/BDNGQ1Ko
M9ebPgGc6dJVqiqb7dBqIivqQ5+La6UwCw6GN5hDBMIHcqsTJ0Zbjs1t7ZKLYAlGT3QeGBmYZG6n
KN5m8pHyMf+P5QtTUyGKScYjx6MenNMJQd6slLpDFZ4QDNFZ39ibiTR4+oQxEHzQPFSRZoXfGdzE
woiF6ziD9R0FeRkf+DogyQgLWX6crRy2HcYEm/+TTICJVZZa6pdhQXPd2jA1ewK2jv7UxBF909fN
M14pHJ9ioSOX0//4C9RpGmTka12quUIZZJijWKsEMqPbwj/pvVOWZ6Kul5YRyyrR0jZd8LIPIt1A
MJFYBkCF+E+R3igafSpIFiAeyjM9WBlN2US08PzX00lYj/enquP8ivAbJg2mkLwxFKESbdnRumgy
cVqWXTiZulw2mNTetlo9PM4ZunCM9CXrk/tKGausiXrd2e7UsUFkWIJQGMlWJ9BnBJ79BcknX8Pw
jC/yxjaI9vFgZv25fbh4E7/VKcF76lgmr6eRYQAtzFvp4VVJW2tQ1mZMwWT79gUULkZ7W6uGYh2y
LlHownUvtF7Kgs9CvNl23bXRucS7oVRu+32r0bUhjqiOCqCcl4wAjOrM+VYMS/dSCBwVaRdh8wJL
k2GgaMFkJt5pJXV0qHu0yolBT0LAjSFtw7rMGAxOPETKxGVQiLjY8W8aQgZTNepyHrBhhd6DORvb
b8Ti8udjzaDKCb561ZAnRsXL4w6mcmyZycZH9xbD07Oix3Ll/ZoDUmIqM98JMO0HGgCeAcfEy481
bUSkRzxJQwtr1yK2YMuARPumGlojaaSqLhQqUeP5i9CtoE1twpuAcEkZ9d1F5ZndxqzR/wHiQ5qE
/dMTYZHAEe83aiJlrL4KdlFT7jJ6Q3ZnZC+KzGrfcIkLEkxZiuWmsm7vUkw4Y4B2ZsgGS+tpWF5x
K04/cQ5/adb/JFw5zNpbI4QTP7meTUFX7zFW6/jAl2jn7Pdk1o3GZ4/U/0dc9G+XBcpx96Sr908/
8e7iQJfZ2GhQlF+E7XFNIBAMW4onbxx51DuczH/71HzhPzGQQLQXhe+0fslzXOICmjXCtimoYN0y
kQ9IXmxb0hVpz/izGl0Auf7P9xvJFHNHq3TEDhU+SHqdNXICbQuoaEblD4Kwu0bkvgUENRFqutzZ
y8+3QWFBgk87GUgy/Ejo3WOkQS6NTxLETplm+69go1Q8MSvBEHdLxzfiKQigTkyUJUkoviDyA+0v
G8s1zPfoNtYDW6zQyK7fFKHZFNOoztur4B7qG3Dj0elQf/Pwf1lf3T6u+BtMVJ09/TR+GaHey0Bw
3Y22z1EfylMBCc1+qp1/y1ldiesikkitvrKinYcEzGHYRh2IiX2hAPjYmWxPnWR2I5rKYmFT88Sx
4k6/doS1f/Vt74i7bm3CBi04DqFxueh5mZrqov3tayBYAApNoEa+5ZbSWGIxRl4rd9Vq7VObNIAz
APAa1PUK8VeYlFqKHQG9ZnrKo72YIhUxSoiEO5glROg12cRPiwlTwHpiQKcUfjphWgUfonskaDVx
YhsGvMtfhIC1kHiRvduljCM4qCarCpTBAiBiy/gqVUfnpMSn8yRzHSyvcnWQ7ibkgbZPUdorNtRs
STZonjZoz4a8hvIVEN0iP90eDYU5HLJRcL2iEXDSUTFTk1d7BaT7VB01NgNMrfYWaBnsPpfUEXhQ
rxjQDaVsHfyEhwNvNImuiwrCEt7tw/ityupCiX6vAQkQH+1QGQMRpFpQu5OaT5EOupUgjIOosbAz
/pdkcXwpdIOOzSJyb9IkgPeqrpU9l4bHjpGgdHcXM0wOlujjIRNXf1DKBBlvMGLtmKNTMrv0Hl2B
xQFD3SGfmqSYPzPq4Mjv07mcDN4Rhd5fuqsczR3DVY/4zpN3d9VPAz0qeOmC8BDrEHDXYaRhew1z
D3tOG2xkCOwKCy9X0WdoBUirs7sJ3d6xgt6AzLFogz/HCFOpHGgKKKV7UtdhUZbD71OdjG/QjnA2
6rqvh7Jl0Mo7bPnpkcycT606gCwdO2wEb4aGmqE+AsRgKWjqwr5fbjyOx1yFnF89c2eG9B7tPu25
xi0olKJHhevzm9v4LNbPsHH09a7C7c8r1jWVjQDQeoHSk6UP0vAhHWRajvpB8JTXwh3gUv7K7PYh
+JMLp0i6EENRITZHLdSMFHDomPYdPM2hEI2akuztD1389Rrdllq9Wm5Gs8GRrZEqclATRat6ZR/P
qbL0buGZ8t7xkCJ8eZWxcQICB1U17aB4FgLWAJAIp07Fm32ERFbiI7hajXSw8I1PpCenqOa16lft
6HtiKTk22qtB0RJKmRY/mTPPrnpaHdgpjAJBlP3beuXOojZiG+M/wFfr10jcs11vDof+ZG2V8Mt0
xDe/o5Mz+Au+FoUe0OwITMSYm7Shx2/VcqmTqAIDeyMS70pla1GsA8bRQLSnAjwDQO9RPr8wBDxx
ieqrVp1zzCLm+vhdnyPf6edIjTRmORBz+X+wiPWQGuqetXYr4GQxoBynceg8Lp+N7+cT1F9dN9JA
eN2MQPOWkYr7H4MXpqwym6U5NyVckmNNtQlTrf4SAff1670iE46q/s/J/Smhn4GJD2Hv4kz9jkGC
BN+nMNepo1VnYh51u4yw1BTRthZ7Ez0+XLUfqvzW07C5Nm30GF/6m8yrOv7s0te5k3aEMFH++Y0P
5O/FLFcpeL0CapHkPK2AAn2K595Vr61OaviImdaDRgAC7eFjXMbcHXBsoR1+Sbia0lAmW5Iyk1Qx
THdMkpxneK35n5W/hh6oqXmkkWwUr5eCSOcVnElO/BMiEiiBBesgBi7MZBPOhGng4X/5xWfBXrH4
VYGHv8OYj+9Nr3mE4Y7hCa5v8QzzOCtkmKRpEulhuOTsxrQ61DAPNqLGfNCzItVP9rIhN9n4dTv7
VSJlslPJjdW0eWT4Eq7Hg+9Q9DvFHjwo+uYgAD9SlnTJQzmBLgYKMZql6UJeSjs4C6YKBJhSZLbC
DsR6fBlRB4FAAoNKmUBCoQx896JMBIZDzruFVQoiJGpZm5axlaLECEvpPfhG9xNizfdRhuZL/dUJ
wc+EeiHtPThtw6tzRa0HCAoFK2pUCA5mqR+S0sKZaBdXpXRpzKTZdN1+XM+3yDWzFI8A/0gB1Itw
ZQfA1O2mPKytA268bc20VCZmCKphvSOlXC4hMR89VJLCxGqjTAKG1gD6VWMdC8aQQiF3nlav/MJp
5dEwHy3mdp/sJLn2xi4E2oZzndBnydMkIO/slS4neXqH5GkmYxAstkyTVJjbipzIw29clY7tFY5C
kgaOES8v2cS+oPy764uKkyS8TUecLNAsiyEcSFf7vYBX9d77e/0oWviPY5PBcScyBV8vudnCiMUM
0oAt180qi6/nEf8XVmnjDXgTXM41J3udPwRd+WEp4u94ceeje1cfQCV4xr6U106rr5Yv7vH6t6j1
SFKrRnfbMQ9qUcVdOdoORhJHLIh2GjV7ElOKfbaZ0SB0qgb4yqzkiEpZqAXD7wCIBKnhO3vdtcwl
bdnIddrFoxL4jZw9xjmZU6Y6Z4UA9r0NboSTNXR/xF0oMKu6xKRN6bZSvTXqa2UTgHaH5d8iU+aD
nTvGyKBgmlqmPxwovS5xcFHmWBG6T6soX+o0sjnyl2jVlL/4/VWZinrhsqcUyDPkz1D7Y+SwoTol
EmuKNYCn10Xaj4dNLMW+KmBibvpMBmZaccxxMZ64Ig75HGDGC79fvyGfnwgmqd2eCj1nFEcEbo7u
bu03xBUAoGEN7u6P0QiB9CIp8wPjEYY/XW/aBdQtq9zqZboqUxvW1aEFVL3LKixIAsT+WQQU5Mdg
ps+FF3XqYzDwE9co7Snry7U0qEuPGnmQJzH/efxjVpMmr+R2MwZ2OnAAiwcaZ8grSRa7osY7rvTe
xVPinpYf1av0MyKNN9uk/TTXZ47xYy394KujaFxd5OXuOoSMbT6NyMNZR8heHgNV/v9LcoOv8XIC
h3RS4EebnE1QiONK3Y3ykUbESy3xi8cMk0c0HI0nAWJY2VeBdnXrqBcsffe7wpjAu0SjMJfH9u0/
f21AHygUTAwQQpWLkLOhwcmwcOolLdp0F/lPECM0XOGf1bKCNmFHzo56STg79KLK5WevGdBUX6Qv
mY0LFGUtyXyl785MFOg5OFrGdmU2hVfMRJ123lDSUAO3LxNJBvRBuP+IgshGRn+7o7q1uUFtd09o
GWI/Zrt8AnqV/pSQkombmaswgGHKRIyADD+epjN7UuV3i72BcxI4rxDKkdJeEvQz0F4eLGR3Jchn
JUTidHdggEcPvsJ779LsO1M9ZRURCC5etGrLDzBGIaoxmFoxbAhdDW4UCJKs/o0pRgVpm9Eti26C
d7GzLJtq4+AkD74HdDgBaLRcXvHtZoplL1VAVwf/whi4PdW1qN8N2HvlOlXngFidrRJ+uqGm5T1N
uFJ4zlgAqWfQupvrjgazMPLah0xrVpj/ALu+G4SGVMiUkPPvbqGNyMG1rIu/rk07F+7+c8Vc8/Iw
ZvooqglO9t+hlTHKhiILLbVJ4P6oGI7ZkeD/2Gu/mne5DMunLpbLWG4xaPeSJa0pCa+3ekR7J0SC
tD3WyQVNbYBqcKge26yoK53RO5hhy4Gyqgj13wEDsqpNFgp9zWbF4DDPFEil0naf/EKPk69Qs9uC
k3QZxwQMMxL55cXhV/PqvoIvv77CrQEj6qVvwfafIy21YsN9FLtqrxU4tyHzuP++OtEvQPxWFpQE
Lcx7MeapRuz0zTX+IQL9459aZtqSitbftNkj4or41F0Wkr+eI5kMqw+IjG7IIWY6g4BJvEloP16c
3sQ+PWPevMPccc7RlzD5qXUYodaZZT+LfR2pWvFW1gA/tual3M8/oAOgUCxNM1BxoiAMTJucRFTa
jpYpUsmskQyal612R/ykNwV8tvpv1O2Rg5yAUV+eSb/n/hWqLj7aMGfCTIpzq1st86GnMrZsVT8W
QPaqG0obL7XFWgMyISk0OHcJXlEuqqlgi+KG9yDRMM23EzGc0lj0sxFD2z4XmJ9GuXhBG5hkJa+A
QG1LNoFVEr3H2WhTW3GGAswyUHwFH8OpBM9f7bEEVbNm4DpAP69NiIB4KVbkbAB+K2YN/bGEp9U+
bSbGnM45BQr2hYlfutFA+LKnt7IW1pVPxrrX8B6LoBpFp29I8k1X+OHqbvgDwEFlvfFHswYUF7il
6EMy9P9GQpSm+HepOTH+x/SC0jToRWqy0pA7ykWFTzucL7RO4rSTA9KrvAKP8J5ce9Z9ZL8g7/7d
K1eKsaodk3DzvsRCkI1ki58bInj3h+SotVJniYDJTczV7M8TUmETrNHh2qmpXhtM4L+6S3xePvQ7
jO7Eb2TSCRviRh9WKGMXZzMwNAZrTW4TOt8qq0jgDLFnt1s34C3m46IY1bTw3cEeh8mfRTp+Dek8
R08+NTJCpqFnY7RaRSjzea47AknnZpw4wThPk24d1cOszzhf27cmPaEBj/I57EHepxvoo0k+aQux
zLLMnKU0KxX/JfipJcntfTZqI5cYu39u+4sWcXP7/5EIv/WpoKo6niDVEiiHVtxLNl7H57v98T5v
GP40jqhO8BL7aw0di2ECa6UMdRT15tP3U26UIMJlQXh7Jpn11L831TGGNb5UCFt/LM0XP/4Ibya9
QE1rTSwpHx/82JyYnk2z1IBp6l03A5xePvXGU2mzbsjDqI+wBSUpHWjCHTvFG911092ERm4qqWbG
OoIfHFle+JixPi2BRfA8am6SJbbCcD9VHetwp4wh8QNKifkv/pkm8aybT6v9a1RmlITjh4alzi3e
n58srLImuEX42+CNls244O3L54EwYKlqtfIPjpj4bz5oTEZODNv/K8HaXDnZDCPcAuVC6mG+7ajS
C/pFkkYo6wVMXmtayXAGFzV+TQx9JScI7p5Pd3iMvurR+KOSf6Gpa2nr7wgxd8hmV1p8SLAjGYWp
KwIVbvGK2YpCGKBG6OYJEurorT23Riqa7LPv7JXcKuJjgOtXCy8i4pkLFXJ5hnZJ/nHsxC0ILkoK
clUjdNvHMkKaQstOxKIZpKkJWY2CBecJ/eNHLqjWdivXVT+13Bt+nAvc5siYBPITNbM8m6iL5Fve
lrwHJkiNsRpy9reE/gXCk4hcQYbXPJezxxu9SVMkhM9+4cMcLxekpdnk2ZrrLzEn2mdUVj1IrzGG
okB6nwcGvIe/7lMstyfAI2xmS9pQPGEO7nbPVG/exNX+P/cm5JpjiXG60pu1bF3ChwNCaBtUZb+D
4RqDtTZWVKwBFsgAsHOVmzsy0G3KkEgtjEGuePcLwDKNgpSy7Ig9mHPHm5cJS0pA8dqNicAO84O+
2/lSKfsBiFeeGJztRWgg1RlBfvdFtzjCSlEwYfqShcNywftczNFwI0FVQUoJDVo8Cn5gfjpsZp9N
dnO1ujPX6y4wHqDJec4Ufud+hl5a1rvGx+m4ahLraEdyqdLD9AEEwcltTKFa4PNkpmF7SQjY5QjC
mExbHa3Rmqzf0p/C83SVXiGoFYJ06P8LAcbRftSWdMxjAU5nB7QPfCkL9iZIvJ2S1FVxGywMcjKQ
RjRWrWncuYIOVBW5JtrL3D3bOS79GfMUBLRb2VsB1GkkG+SYB/yzz2moK7SbxnjZjbctugI1yWaw
XtZR8kpF7jfTES+WCQrz2alBjUR5WSGhlm3L1Oy5OXTSBW8qHOatlnz4WgnnFz+JdscRF0enfwtz
wira9fh7lZOMLA//AcQ5ziTvdS1UjPDVDI/aVZXGyEE0IawoyvC0nG8sCnSBiBHbUqINxcAaWWGw
gwYoP5RmSz6ng+/1of0ZTa6gTUVYwyseTd81g6I+UAemV2wlnC24WKMK/Oh6lTcy5JFBYDRZNk6C
iJ/LBvwaYPohuzY9w5kPr1ut+8+1xvwsHzvwiLY5n7bFftn8n9OFCVx9ZsOungbP+zlVJp2emXm5
vYCh4QdLxZqcUFMIUAssmf/hXLtdi/4klIvj3f3XPpkp7aygx4tp7WwuOu5E4k3u1Hh09YaOv1lU
WSImSlMEBgcsFWjEAN3r9WgD9zLOnRcrvkBqUUZSW/KsCchGSNUS60PkWLURK82ynRP5yRyWPgDd
JVRFSvvcFpK48SEulCNDtCgMWFbFd7LyNEBT+/XAbFTslvgZ74hENVqXvQc3iwr7Sc7v25wE63kF
vMhrUDZmN+BY/KdCdrjXHcBZtdB/m/0x1osi7uLWQD/giyETDqiBs9n2jevkkJytCUTNsGleERfq
gUpkDrvsQDSY52qW7kjUuO/62bWBC7P9+C4dZpJR82t6ptzgn1X+giqo7MJOMojfwt1ruU1qG3ts
/b/MlGBydD1kzDT02UQqpzR+mABj+GormgG7Mttha93ZuqhVk5a1KMesjBB+Ewkn81guSA6fRnlz
bpnreXzaZw2G9JAeI5i6DCnxzr1ELkY5pE3H074XCeznx4Fda526r8ktrtJ+O5uYmPdBU1EhpN3B
NTaRgK6c8e5tcM8p84Gm5oArh5rq/bKvb3W1JArahHznTwLdS7XL3G6qhwhIGqk9PZRWC2Vw3d7Z
OaZB9aD6R/UzIyjX0S3nECHlwUhroFS2922EcJ56/YDX12qr3QU8CxFkNGdqLma2Epj9WrUWovqJ
uDQtKoyQ1V0l6iH5aHVi9ZN7vDEXwDMcmbXeg0zzJOuVtXn6n2ubwq5aBZTvELEaPK3YmRMMwknM
/m7G6O4rWyzauKCu5CYSM8FO6x0wTR2OEMgBy2EgjIJ0A7Oz5xtTg6DhWabeG9e5vJVupeV7b6eT
PNlwE1Y4E9t00dRW9C7y+8hJ8J+ckBQ5vU4Gh4jPXtONleSQsI+ytblQq6lxIEss7Xesi2c/vNd0
ET9oC9fgf2aoAnmUEGQoFCx+fv9mOxwM7CE5FSVGjJddsPriYnHNbLhzZevca8vHv3GzYQiqb7Vb
Cd1ualRAEcUpD2uK1g2q+fEUb2KbvOqYRGcZDae/Gf2G59KDJ0LvVPnezzmJaTOJZNNRZckJpU1y
57aRixp+IRkxSKTaR1STzSI+46ylx6D4v5FDC6Xc7jFQNkBnJU3Fa1R/2K0GEK4yhh27EZT0qwc4
ly5O29f0BBuc24SNQoMLdoh8UY6t1hg7aFHYh2t8c65GALsQ49H5FWQQHwrwS9ixBw//vHpgSVgt
17n+ksGeKrM3ux230QnaiQOY6UU4vFXfNaU9gTdtKeP8B1JuWkU+nvWnsAhmQXvHp3sp/oE8QByd
VoD0yif+0IHOYMXNRNPm7IJXqMiHVT8TANUebO0641t6fDd/CUQJKnUrvaPVQu3rP58nP3u2zNpH
/H+mJEcuVPXi4tgt0InuR0/08XCnCIzhk8by9mU9dFLfbuA/G2UY6Xxjyj6kuN1nK412rC937N5v
kYAxpykAziRKRk49ePNgQz9kL1IVLmZe+XG826gxHaPo0J0hG7w0C9Tqu9LLIdkN5d25aPHiDQio
QXLwlBPiWoqH492WRxWvhGrSjLtoNlzwIJ5z8XevJ0xdYzHyfInwxpIr2q+O7HF5/mYsq03QnMjw
3798rQcIwFoSxwwcHD/8M3eFPUgnSBcN42h6m79LYzT5vmq2dUyt6nBUf7G4aa+MMg5lzbDwk+Sb
PZoqzFhPT94nVjvJKzYgpf/AC7kkMqnTxGBkB990x5KWKjhKH8yTWssX+Wtk2LWlHyVYYfWy9Hyn
8HPoasljFuJAbYYbH2HxhdJ7TSTX9pJFEczopZM9/yaCGWOjFEhyfFwlSvsArZVvYwGu7RJmuBUp
328FJ8DZY6UM9VW5IjuckgA+MmVvehhrnFaXDcGqdIlrNjB8rhkUobQR10y6ovg2py7A77latja9
dVy4or1Qxx2Wfzbz+stRxrEucKYOAau+CtJrNVk95e4Zf8PWqu1/tHjWv9iO3FsLaJ9Poq487eSU
MSkp9N2dC/3krmCPFTDEQhmegKxaNtAmDb5Unlp9IqbT8J+UZDDMav7VAr7rkOfxyTw7PNt/M2Ip
vPtB2xJ9z37FYNlKWQRL1bNd/A1Sq1Tfi3is1HXU0TVKk+uzsoUq+lVhS2WGH/B1iCeF4s6DttsV
J3DQjg70C1sZLItdZgSMZJP/LPPolEL4em1WcoqZY4MswF8/Bc6FwSHxO/q23Vfh4CPPmRGqQRwZ
2Q4Yp7anfiejVOdZQQoHcDKhi+fY64eSH0OFI0jLPu2Qm2YeR9SxzVreYWs1JNf/MRI8aebN9NfU
bznnRjux9Z9RQCLmOTl7aG6LLjhRFQZvZU26SJIuij2/Z5dteikmSYHtVgvc+lwkEax1tiDPfCLb
XpnSNi4Tr03Td09Oe9TlfwrqasHHiA0GexRdcZGFvDhW+7okpSwa7e/qyCt2P2iytFRK5lOYcsiS
Rlxx0OH7B3DaHxP+CRwLKFQCB4ciSZciHODBQ7mHNi0hctoABC1odt1S6uM3OceGklbOZ+og/F+L
H8IGg2l27f/El2rJucaTCn0Pdsuv6/uF/qOSrNPGJa5hgil1sIAKOecXtKElQQDtYgmwCcE+4SQY
rt3cgK0PKtRNAA3HAuSckpVu/UGGi2wXYOAaqw81GM5Tdz2F4KrFcy6uz0wk4cH5DCyZioMIeJJE
MxhHLvqPIeMFBB7rcKoEFuUKP0Z0rLxt4yOHN/9D2lF6rf6UsVp2MyxhWOmFw+k3cK+r6KKyHkEU
D/QxYQqDkHnxuT51gzmvS4v68U/WkaT4nggXGS+LseTuyUi5G2Tyo6oDW8fL0BrJliLd2fOCq/Z9
Zsooj76UlqxArLt+tPmaRmfcbhi6262zVa84jzLvosj9x9W36OtS6SeZuZGd2EcTu/4FyXP5vZ4Z
L0POH4OcfnDxK0vBlMMhBNISOxje+P+ilQ8KNIEV5P591s6GV/cIJE1VTVOA30nDZqCd4xkITXp+
wSEn05n4PwKuYOaS5NAlZLOyuHC3B8NlqHUAO+2+sQKxCVHRHm3+e5kaLSlxEL2xy2Rw00mwuWiP
acHfKoNRaVXG24y+YfnAww1c0fcKafy4t8giR3Cv5O4qBn6NHnwNDKaNNtnQMW0IDcH6qkEZV3cW
r55kbgbiPLd8dPjciiA1X59WZGJ55LIMACh04hlkMYIQLxYraQP/WdmlIxK7xFodqoxQMpfD2OYs
uC0DBstmQhi4ck+WPo+T7rEv9u10vpqX0hUWCrdw7OMkdRMaSvKB2tBmxX3jAxEqEWD5qWis3GQO
jx3iVlTEa7CH2enr7dO8NRV8jIUWhyWNFeaIeV4B2TEL8ecdW7cAFBFL66YJm6QDHdpd1P20/ld0
mZnxI5gK7+D9OslysyWkhRhrgzMFsTKBMawlQE/7kfVXds+QbVOSDftcCRkC2aBma/UHMDjCCLKC
8q+fsj7P76A1E9JELN8+xSF8akp4XxlQB5OANN5qz/Mrt0zIbWq65MshNGOuqPYFFiDsOe+MAjks
6vYQS5mL/iV3eqAOG+kBZO+Axc50F9G4TGBY4U6h0sm04gfeFiVsRhHB9issO4uxa4SCvu+LDxNK
r9JGSG6yVYddAiJW3q6VTodRGP+uIDxBpX1e3hpWpoBL2xerlcqWJUDj8JxQUJKuVtlW5jVAC2FE
YRn1EIULwSNigN20aQaKHxKiqH7QWswl59a4JLm5sayPrsUlPVrAZVOHGFMcC85sHDu0PcpM33Fo
Za+gKSRV4M+TpVfFVeYnbNMWcFzUVnKldYoxRQ1cLvcSQwVWc+/NIJoSbl06KFKHBbrKdTDabSs6
Ldg6TtKIc4elxsPxvh7y/9jqw91UlGe6Td9+a8XFSAWwWsc4yxWnfSLFYuX2tOxnmsmsXuu4RaSw
nag9FkVhFqh6BBi5MzQkDGyjreqRxEGfWLEIwoSvtljwBFfFVpQZneBH2AmhdXqVp8uSMba5OEzL
OXZYwPik/nVUt9xtRYBRvA9LPsGC/3JsedvGZcJWZmqEi6CM9Vonpi/yNPTTEKQ20rESgy7SwzBz
5fEDdf8EydTjEFTkbE3CaRt2IPvCS8ivedPsW/MhsJtFXz4KF08e9diuG8BXzup+kuYXjSmoI1hz
p7O4nFFPwr7pWyMVCHgRfXhtzPs2ZDakCmXjlbd7lGcA+visOxorSK7JDvo48xIamEbicyM8P69I
tE7mUoQmGCGmI+dpHtyXY0ROXBibxElnay4JPzDAaIM5P9ewKQ4DOC/yYHWXAPtFzumLvacqcB2c
xK+9QIBYVmCv7LwzhfxTFx06rTbiKuZ0MkRUOAiMbRXOn/TJbrkXoFv0vtEVfQ6VTb+hVvgZg+fZ
pscKEHeR76OHSLG0GNQ1zrUQPdOi2mlW4GldwZimJSZeuUqP3kFlPwrdNOE5gfYQJv/xtkwGMYc/
8MTtK6KPMe2H+DyozLjrrFx9CfET+T4kgzihZi3OUov/FJhXCsS4WvuS+1AIJkfYzHNy28wpfb7z
Uc1i22IgmO8G/RGMmWW4ql2YI2MYGr85qdcBSSD5gloW1wd38xb/ILOKKSArvw9vJkTtWtQHjFC+
lWFreGfOLqx+/G9gVVawZLXfqcRvo1tOsA+mcuiHjS/jZnzUIPPe5f/cR9BVEaEIk3yIZMl4Fgzx
vvjJxwmbiqYwZRjst0GrqOue0R7CRt550FeCeMTTPDjEZHtEkDs4vpI9eJFnKHoODHyJ0MP79AG9
Ek3jbFkSMCHJfmXrKs3IUGoSFkT4HWz6IUUM9IDuDoeJcISOF3vgpiXg8DUBN8mvz9LwTTij85US
dpBEIKr04Ve2wApFcd+A7ox+vvmE87Wb0yshT+RD0M1lo4t6B+9TCa92AONiLLwBTJEU6ebp8DOP
EbDTOdde++2in6yuhkvUcJd4erjLpcc/Sw9OBNhhZFPWx7C21QTLOxBFC1hdrc8F9in+1YLVWuH0
DK9Cu6P0X/Lkd58uC/K5OQqyluLU5HdsBoImpEt7Cw3Py60CZ8a+TBnXC6hcelt7j/sJuPPGLSPm
dE+mrSo+3zyro2lECqszBkc30Eqg8nvSfRusVeK7UlvPD1uUPQwIHhh3uyCXkrOltqefz8z1nZsb
DhYtv1F1k1/ij6oU4r8HpGZHhVi5CETwiWbsE2SXR1uRJmDxS6ULULV9YtF4I9gPYDJ1wnjj3vvD
bpkChXjQw1O3ZvuKzuyobTPQiMwOZgc186dz/rimMsHBW90AI74WVzP3iXSXUBGQ55KjtOv5GVpg
Ny7lRNTYlC+uxtG5oZj1wsIfwh8rp0uNdFAbnZ7XiMGRceBe16aS7z2/S3LZUgwSM3G2x1LP+T8s
drx27NjADkAINPo2c4anIzXvhhOFoTh92KpDZ+aUuOwNNDCk+CPemZa82DosodhPbTrJj1ZXAIdc
mjYjyNYavwWhg1I2fs6xyr6MPr2+qDeEP2ttPXWyLZIgZOFNj7fdaihfeWIMKJxp5c88YPebUYXM
3CbL1ZRGmEvcGdJe+jJm0XbHCslWGrGb6Ykxs05z7HoPc432AHg/dFkVD8u79KpyNZkF1aJwjpK3
THVN7goi/OMT3Yj9SYDpypD/JWMH5bk5G2xNiKju1bs6ka2J+LRnoghfe6dQagpRnVn7DMdNdVn6
OOCJZ5PPcDgOfUSMJw05yyT49zfUGu9+kxMnOdHrqEINiTBeygNBn97jKd9MoK+e+U7HEXElZNq9
dYt7AMwGVrWOKdfuAhV03TdE3q4Vy+kKurYR57LOY9768Z5UAr08sIR+o7qbgLi/gAT6DjQhHz0S
JtmrUmjn6LL7INoaZgbmaAr7GxiEX77CvW4st3TV9fCHJ5pgcWzRuRpxCn7kjOvEcD8T6d4SMEJK
Pe8UDihoHuX3aa5YFoAkWFoTldoOLT8ekWYey2vSqX/DkUim1jinqLstLZi06DSFmV24TIGqeHtU
W2/f1A/kyKzU2zNP6ZIDI9qfXydZ1n3NaVIkHsfh2YE/xUm7jjRUreR7qOHV8RAMLj1EuRsiKTqW
wFtPp7wtAuhOqmCoL1OMYcUg8lgtWTs2OySdBDmd1jHFGnz8oCzxru2moZZT4MWkI7K1Ab8TI4YS
N6hBs/Ce6cXFIaKzaIj2xpoR5IPoHe6C4DhkC2ktlWvK7qIYbM0G6reRrcWWwjJH2b1hbuIdlHDa
QyPvV0meezx4w1Ri/cUFl6xs08cFtPtTxCz/uswabE/XPR0iCJKqfXzJED+Fp5b8qX64p/W5hciK
cjEIgm9FNGnV/btczpkZXSvKj5bv+sLf1ZQ0ImHS6GgxntNtO+OGyRzzXO6GBnZdX/tn7Cd49nJQ
P7e03Q5ClKaUMryW2W6LJumvKk4TPy9xyzrMYG3AgXTFG1IsCEruzsg2ZeCOAd6N5XYbh0Fc3iP7
V2hBPXDPo5JxeUVDnyOHnYdpkd1J9uXYrrvExl8ozxnFuOmgm8WJdfLYAxRVstDE0oKviwvYS8yL
uM8xv6EACwCrtvKV/1f4uU9/YhzYEk10duHiWCwmivH1VrsGC4Sw2wG14qPkQSplNa42v5vB4+m9
FCziaen224hNUdhjpsdV7AcGYwTVNEy/8drurlfDgYIYHf48hjHuLG4bp8Qgp8AsNQcrnVTacs2i
tOCle8HPMMu+z3fY0BrXNpHAh4KGNSdAsbr2OBkukw7t/59T0tcN7OUd5eMhA9OuDw7cHEpk7ROp
ti7zxaS031qeHRBxw0dPO7EJV0nq6gNbH1KARKV3k7JnzgiPZjjx3DWCg9yNyXBhNxIIkqs3RyJw
G29lVpAWgkWEpgjZzn3xZSIPTU+Kko0yVTcvL+pCKZYkmr5ujrWir3SgGPwCJLnxAQmgeYeWkkZ3
aFsNwzdC2C+ZP9/+hJvVMPJ2LpqTgrsQF7XPMLaGUV5TVXTWX0/JmVd9CC6rpUcvMcP83kWOnWTj
qmiyFe8WF3YOUUAIqdcJ+aRTZs5tA1bw1l/3SOf27pvRr5Cka8XAs2fSCWFQ/oJMt0eWuyIYlILT
6SNEVTNom1u9562F8gQw3jBpm0zDpsXrZUOSEJBdLBrBOOQbT0cXMlKQ/rkxYkg2+H4sGPLtrStL
BuojhyKPNKiPhpM1eyGinsKt/7xZoNMCCzpQvTi1srjz2ocQP5r0J/fkhpHgokX6WBKRgAyHO+Tp
0atY9BiMn3TObV9NnfbxahfTF3gIOusW1AyOApM/oJxgYH6jnsIploM30BkLNW8dVAeXf6pk9P2s
dIwxx3JTzivRKLssM7BJn71289WMkXFZsfwWL4PF5bd7c0b9UhTOTbOnaay3RXA6ZwLuWnSYzbzq
jdUPk25AcdJuAjEa9ZaszQHH/hh4Hnm/w8UtK85LUSFPXfYhpbbE3l/Z9uNxYjyqUxigHo3rb0uI
Mk7swuiAOcCDYI2+YuoNebmA/5loFjp0F7wvO062cLckiwS5cgdVmSbcu2a/ElHExrlA0ylXPYRe
sX65sxSZ06q+5Bg9Z3/UI2lUQwABtTbOpUT1cwpkPRhoXmbN3CI8AYr/ELCdchazKFPhfLIR70FM
ACWBRnHjrn8iMF8ihMvJYD7nU4cGrfta2iocECjmTGERhT5yGTbVZMuESGlCFOhS7dS40EpuCynH
C/racuc5hDHaZdr+rTwzKweaBA0TpUxO1MZ6yeHEBNfYF0LzNdD8FAP8lSJQasODNVXT3esMBs7s
f8q4yP5O13Nwf/kJzJwlczuyr910qg+qzrSoOqLzILE60XwyOj291y4xNHdHw/AkOzaoeJEFkK6A
VxcoJP1pPzC5i9TGWrLgK+P5ciauFitLOZrCWFfeY3i4zvmA0OgPQwoHXTv8jDukbZOKvFe1Bboj
g/uZNQPq4QiYXxuT94uLPGBYozqmZSXVh/KuzMKx2Qjwcgk3pvfllW+rV2A6QRrKoeaFvFpNqnsq
dBoj96Ci/LlHwhQi8l4gdL/HSaen9PHzvmxKmTtsMXYkr6T9ivy6VfZWqQYO9FfqDlLbvAyXwHHg
x3vIQ2xVzx2vVCbzzC3dJ4jdm4ALLMRJnLXitmNTkkKIVNQJD08qo3nXz2BYL8e81ZONTVbD1fhq
hdgxVTbFDVUf6a97uwFNvAHN9l7U3ZNaj/8zP9muAZ4hem3V9MDoE2yNH76vZKKWp56M0+R6+tCK
SR4fMC1sGgBluKitvWmoM6Ra1qqymRbD3lSnSC8BZseDVpG7xgVtjXQrNprs6h9YSghpntGopB3T
R6Qk67r3aNWSXz8mdaFZrm3fKGZKXLinEtz2yCsKTGnADKSU8IZIYVgI5sCi0ix7UJI7mSDcGxHL
kgDpKoFxJyuEmf3DfhtqyTjGxG5m+J6KhNLnIW1dr+wAYB7q7Dd8cW09eVto66N7cs5U733vbFRR
stNdVg8xJ3HQQe158H2GtY3/g/dxPLRVifbizaHF8Nldx3eFHgf28RcOHAOBVKkW6evfMsDN+07+
qjGIMFK5P/2vPoLhl4nOdpvyPaHU+NkHnPRwOOw3O747TANCd7R1W/MtngWIk0zZnhDm+o3H7LBz
YdpKPW5CBiRcX2CdXDzEx7EfLSEj2RJrs4amxd0qHn1C3cgONfRuCtQhYTFc4GHxKLXq+ReoGUN1
rnNtmSpfeJ9K4UdhUiodFhWxMoANIuU39NOS7CY3Fw6yc4Kr1iLyhM9i709yx3V7LOfYx6VyLRHc
PZvfsMM6WfM2arLenbUVDZK4p2jVIQQnUF7kAVfMCaE+xNNJebrbH/ySEcPT8ZyvPswr1aHHnMjE
4A2GFjZO9QKLbGJfrBhPuq/Gl72ecLUkmh9BGWjkN+ruq2aNi5xJ9kKqX7yov7Qqj6Rp/1o3th0F
N9Ie/iDyUA1jCkvaL+bJQSKSr5tMIqFl4cAUcbbjbn7NHq51P6wsD0NbsVwjdklCFOr+yYAIPKzx
itzcAFTM/xjDb310Ur4bIxRln2noZNl0T/h73Ua324cvfU5ickTU3zIKWhuLrC6r8waQZevSolRr
17B9hYxH7otgG1z0Fnhm28TjPGpDe619a8i8PtyiflU7VLFn1t2PImLJy9Ube4PihUMeIOnKfh5r
SVwZ5T8FEScMbMaAXfWcx7IC4aldxYMk2VXNGcdTUzfey8SIJ246qbYjCllqFKDeoaE7oV/btZEW
Psz/OZzpfdzqw1bfCKyw8CMxtIaz4Bkz+bEjv8Ob41V1h0RdlERUspoKrXOMO5BNiGNCLrcQpSd1
iXQpCts0YdK+TTy2gZfWSkg3GDSxYlBBxMQGwp+XHfbRC/CSNSxZV8z6DY+EdZ46IWaEGWUR5Bk/
tOoOKwT/ORcxXRK/EDrvALbBJnrVCCo+OyvMCAlCREPrAp5O3bxFZRRBSsNFhxqpbT8JM7iAkajz
GI0ZFiTfICuC0kkhjJzFF2na8zRc7C01V7azznq0zvAwlBKL6d7fa+ndM1nYbi+903ptLv0BgdeZ
hlmVhAKZrH5qfSptbworRU61SU8NZ5jz0RIpFuZq8iCsZ38FUaUiDKk5ulJeqN72yG80i6KE0FVA
qigXhdf846l9c7Rl/YYae/CfHJw9jLsXpEmOXIZ8u3Pq7XXaCxmiEJp31CeFh96UN4Z7Vq8DbZzj
ohRVNanuual+OFjMQ4PFudCj02RolPeP9BCmqPEoO9O84Be3+PHRls1NbKGixjhJe7EA12KyZHFp
pN0EB03NU+Kodnz30QJsognIiBHVoL3gtZU24aslFL7CWs8NAVQFqcOwt2Ya1z0XiJmnq3glmMUS
y8GarEKtoTbCaUZnbx5fiCGyrWERxmeiJKnZpB+iLZBmm4lL2hUReklo3gtLF5vLaEFH6rQK9kZb
16YTkLFYWyxXL/kIRmJnpTg6DHXByzvqVQR52f9j9Qg2R4UqOVPy1F4U3svLYBwrRk3yH10GgkEV
/QXU4H4BFKG0fMR8VZ5V9vmBMgMTp0by9iqgXLtKRwE+Vi0T6o0WTgRV1bEgjOiec08XAZfeoUSK
zhysPVu9FiCCk+EkoDx/QGH2iKWetec9mePfaNLELBtzzOKjrMwzzAr+LA5TjMcoROHV1YRvwGPB
yOyIMJ1ybI6NZNhnqYz171s4bs6LZeNsIZ8gtbGXyi3dvWZuee1PbIdaRGNj6tttX8+D+GTxUsM8
NwJToO0Ak+6Z0ZgZk3jE17Sh1fHb2+zdRaCB8cVjt6XhN72NYzGj/7ngyoUykEeZLPvBzb6i5+dE
X89+xcaQWq1ab58AcNnON21txrfuWUdY7cWvl3DcTncxjlY7VKz/z0p+YGzFLHqKeErQ1O7ELAAv
imcN4vcrqlVcgZBe0+Jo+cR2dCPwmuy3A9bEhq/32kGcus9oGiK6+IT9ccexS2U4xbv7JwfLWpnV
i+BFsNFvaTZ3Hf+KaBAqa3OXoBgRi5pW1GLs7jnGuiXcDdhUytD2h8KWcHedH/lKDTggkYhPq3jH
MFPKh7wpA7yUmwEvM4VZBGPMqLXSffOBuM2cWYQDDt0Hc5/mAKEihnI4YLhrJzJPFlW6ikSSVPfJ
29vcfCELqdEYc6FuBKqxO9cgqnadG/b4BKXbFS0b6WYgorcBiQW7+UhlejWnBqEwgBu8x2Su/q1Z
vT0F4px+fOieiYkCVql2MsKH+Cuk5W+C/arwWRsYhzQGVvumW/jV68MlSDEd5UC9w3e0hh+sgH5u
xS04RhIgqmrcGI4ffvA7k8HJLvY3gONLyoq/+MFuVYPBZ21yanU+/2HKchRK4++JpVJGZFNvgZhl
+KIKRwjWDorZWCBsCfHH7l3gq8dPBk5UqYtW6sOQshqLQtO7ULGXRN88k07+3Gns+vwxoPbz54E4
v3wPYyNovnwayqwgDPe3Y/ZE1NSfOlSa7UStaXkUQJPOHnikXSj5mITK6UMPbgH4o+AbNDb0pJla
zrety801CycSZS9j1mBgKLJ0gKWq6N9NbuUX/DxC6D00MBQ5lPyZgwJCTt6Hf0f3IU4qShntlHMr
EjfBnUaQMl/wtHL/9oCNZk1vxYOmwHvN5w+2eRjLi2jDXWsI5K2lP+qkxWDSSbRP+75mkrbzK4ui
i3jZ4gBj6Fxbl49WD+jMFii8oVinP5IIZKgjZjfBA6ssiy6gaGAHJnWtLKLY+n6BDlceXkydywDR
Tjx+d2/zj5toqG1EBxcdMUFGbyAnyWO1xNmOji7Zv5KrtKZh3JIiDUwH1eMVfq/J6lmoZX4WIDuG
PdbEAHhAf8sjtjec0FHXxrPfOCee35TFIkVSt9XjLZgxAVv1gKeEkUL3O2CF06cGq9gc4Be8hOaa
bPibkHIcTBWoSb/OUiN2Lg+TUVLDo/CHsIt/zpfVRHQu2HE69dY/lgmHtnH+9+a7OU+PNdRJ9Vdl
o4cWmjLAW24DcsAnvGPf8Liojxi1HYd7/o+O+Hy3gQH7uPQRma624MxEmfjeRrJHqfzqbs38CEpQ
J3pEzyFmhrnrDQrYrVIK2KFYOGt39JvSpCMb3/IiE+lRwT08lQuplfzHi7ZRZMN5bC5DFVkXNKXm
xfvhITpJND3Nz3VRtdh6AS8b2RjPSc6zEha7EcFKEv6fcl54xUvcz8oLTJwLK1fMY4kUwRdTWJ4W
AwhfofWpOyoOnNDHAUimec3kdsMLHZel9fWGgoJYRXsqRFVEtxj4KiCE7WdHsIjHAwkXogIksYgj
wuT+LwNv/BbwW9gkF3+sDMxShNmgdoXM2Jf1W9J88s35ExHz0afY7NJurQPi7d+vFMHZ1ui7KvI6
EXLu6XxwHbM2uDMjHwjyrrEbEYP3PE6ot/flPjgDAoIVT419krS5+6fetS5KO3hFP98ZU0LyFiCE
8oUIIHORlBZ3GMivHOUt62PgPUQ6fNfOw84rzclYQ/loYJ+Q2x3j03lojB/58k9P52odJzpblvqW
6Nv7Us9ytLRmx/vtHyw15r18c2LaQN9HpWJ69l7IjHqkpJRtsq2YQ9lsKLUOFzC9NWFZuJQMtt+9
AbS6VgRomYk8m1vnKjBPSVU8brWfMHIQiBr6EhMWPAjxry4SEzcoNwAERZxp1uw9zLaLIdYEh/Hs
rS7wb6JooUEGoAcvjF4wO663qZaHQ5Ao1mJVyjq98YIqtkIC/HD/hNj2KQf2lw9HovYTEgOaBShs
ZGgNlTSHMYY4rMl9LVIDDz6PXsgBz431kBiS+WjrCYrdYjWeghuTHcwDIuGVH48C4IbrF8ZwunMa
CqqzW8KtEDlrsUus+C5aRj9JgHYPHiVRVe14sRtYrhgQJnTEtZHq7Odk5l5hF7OuUb3/7uybzJde
iU7pzsrq5HJkdSFRyjVVmFiT3bw9JhcBd7TkMW0QDOcqWqpGlYC4bkaPEmetcDasTmospNU0uEqB
uHlZqLR3dg3J40QpC12pofRN9F4UxqGgGs1kgQGH0lra1djtd+6iJrkrLqEX2QxLXE+z51umEAGh
OY+qAv71pc2PnBsHaUFxwiTl+hVKfT4qEITZAtraapv3YX2Yn7S+b2hDSmwU+fHpSSR7IBlFSOkc
CIwBpzonJELShioV45aIc945cwPij7vKqaTMAOJavuKaYZ6U8Tw8t4QxbhI/DLKURmVdU6EG/u6C
8UruLRlbX5ZrGxp2JgqpVL1wdFC5WrnWfw94wooVdc7PpTvxJs1qZJdkkswFTU2Oz0Ksaeyc3AVx
Hpv+Mn3yGMr0nPbA2F7f+RUH0bzZtLjDQH3ROQAbP6Hn3ffe4AItWWFClanqvtBqOkEpLLtzI1BT
CqjHsCkinjKr5iT9UdP+qQUm+myvQ3JYrf1QNE89IQ9uD2ahxkgS8WSzvGzlYCBtn1u6GuGOSvP+
4VCf5dHt0Wn/nhA+ccuI01fUqOfLklTsOWkLFaNyX25I8lznCHc/uP4CQ+DuIGNkStaDnxgpd2aG
yAhSBYuh19Lm9YUJVsRZrTvF4zEkII6TVk9qG+xWIb+GuTFiqzuJcCFw3mfT4XKb/dN6jhcFIvL/
U6q9ALzEY9ACU+WpwFj2m87L6CUgmUenfmlcOVLREmkn8lhhhZ0Orzgo+Wt98LGoBMu35MTZmNsr
9IkrE7fgZr70TbFJa8l1zUbZhN78jk4J3Wp2ZO9B0Qmdh+qWOqwjeEM9THyDKjJM1gKl2I6/8dQw
lMlbzo27oxUfQAmJeMmIQsKkXDWsUdYcYF2Hw7XBYeMqQddvoPpuX4bXT8R3mOJlqlewbSPaS8dQ
ITNLJIYHjheEsSsB8SQTat2nMLauP6qENUiHfQNl9uFHSM2zYAn0rChguuFg9dBsor2sD0BFFx16
oJw9r3q/OeCFkKLuzsUgvYJcqS+WjWNojI2cV65bFSEPlTIvTYmcnwGL5hyGD/pHlO9mrBlcTm5K
X8boyeE65IkmvmoJiK2lhaYXZeGwkPpWkdfPuNXzJMRhs1+TU9f0HuVkd5Xgc+tp8tH2a3EOswbB
Q/c6sMiZ6tDDD2PoN471mSsieCS9xg+H2LurzGisIzF0yTg0hvv1p71DQyQTaNA7jN490ynDD0HR
OeTRN7In9HQO6oeFteUIBJvt4x6r7or/Gw3diGz6nYb71M2VxWYrPPoZleGIwT8lbpQC3Q7dXpvc
B1x9ewGDt9sGjFfQ8+RMbRpSWDzQn/QzqkrmcGHE9L33Ygt3xx6t28P2xfscgaPU2jU/lK561BK0
0nmkETT3V9fHt9Bzac7NxBanFmW2frIJKZ6i5W1iZaji45Cq6LSc5/4RiTomFpDUjyIp9sYvlAWp
u3wh6cP+HEmSJq8xOvufrnV6vfs+QPdXGk6i43RttyifEagQasFTr5YsqvmyBEWOmgsqcYIrdTlw
596qiC1TebS02siJyUM+kfwaIKDg/dWtfLyXI4hqvVqTHP6sqkI1O2c5z5SOd/8D+TlMYPtoErgo
h7kR8H+ukLDxcdF51ahxew5PQ1M+WX94WBPduYH/kzesl1IQW8zhOKEdmUMP9UhFRVdA+LRnvjRC
XNdfEpe/C46weactIk7pSvMsdhXd4ZQYx1mjtO1NlHBkaJKCzkvvDPI4YA0rDpKN+GL0g+NhffUH
DDvleHXYOQGzdsdcH0roy3RfdIzZmF3Y6NfRPGnYA/j9YwbxbQVoFOGoL2IlLCNRcfiq4lfFcnOq
R3f7XQPiozMbcN+gZhUy9NElUEGjku/KCaaW80dUFLUIM6aEHqxxxud+K/MZ4UM1XgKE7LBnA+T5
PsOaxWYfdvgz9WE1nHO8UjLSAOAf+A9Vv04891YjngOeY4h9hPEAaFw3C3QGaWUCva7NRXEykeMC
aFkoRY19pBSuIPCJnsc7avYgihtQpyu6Vft2waCXzqNMyDvd85gwKSjG/qGeQp0N3Q16ITAdcutL
JjQJr6zqOCSzdTsyNyxhibreWjY+ZKUu1EyoAJFSqkRoLBiTNB1gvoV1X7ZvRlPI8p9YVaD3Kkpu
KSTVm2JcCxOkKhb0RRqg2rPc+fTl3Fn8RtUu0B5LSvy5IYaUnyRhy7xle+MBWt/18taH67zsU1Kx
tQgtHBT5GwXwCEA3fI2ByU1CMnaEnsKJxCzTo2KzZqHTRUEcirKRkOOGMK8tDUJTPLzgPAPlojni
pjMrQN7RxPwuK6TiqNo6rhkSfJLVduLcAB6wws0GhYrmxwZG86eIAFRhaSFNQ71KUlwPp7Zhfqwi
hArOYyRvaKt2TEl23BAC6QTOPocYIeBc19ZhAj46TvYvJCJMB5GRcLS1meqLHj7EQrvHRp4Z0/xW
OJDHYhbPqZFiV80R9xJ1GSL1EsDVEw6SseMZrut7oVL26cWXOKum30ckvWiQtFzIiEoD+0eKaaca
I3lm4RNYTZqzk35ogMCfk7QT1XBhTXOxZuiLr03828U/DDk5/ecv+3pIfF0TXlXT5jAgCSxjMuIF
kTDEccEunglblP1tOeOT3NoD0F3IfeSRUpTIH2cDIocK7L6n7JY6i3wyjF1yOfDDnO2k3axmziPx
iEu8r6Bm5ae57GtL0ki3hJY1j1gbSNvZJWUqBEs671H+oYm+c+yQoEswuxwEkI4dRWeCQa7DYVaO
PdVScD9IpH5pN82zK6vh9LTWshS4vIWZNZGZXnkWoRizS8XvwomwuURff8maqcCx1ab2B0+yb43u
TI6zVhMviKidOvaAUvkDia0S9ofA69qos3y3KttzTRRGBKIKPd6niCxh+lqNrD13qF72QOWiLsnR
J8GHZ7nwS3uVB7aHYrk/uphsp5HAcjIDevMDbdoRB9P7T9iJ8wNaWnMSaGxdyIIHwursp0f2I7xS
yR6A4TWQtHRLBtpq9sqhe2jYSyQQVrwgIzMFRsl+76/tqHRo9qsGfFJsttJk2D4uSFrRwm4YbQp9
3JfUBghecLwCYFz9fsEL/70N/n9nCEJmm7D0ncx5YHg14UC6VicVA1+kjEOjZ+MVIWl6wLUPYcmw
6E/ZE6FT3wCrauoS2g/fkuIIOLyg4B0ULlcosHEhNtR45zsXpL5hX85hYTq/+gleM7Rh0NRtA5og
UNj4eQoBTM8RRrrJy23M/YmFj+PR+c4rJ/lSFhfhQMdTji8Ql2AKOAGLA1T5yJTSTbQ6EB+k8wv1
FXYUo7lmYrJYtU38cIQ4cDUDRuIBI93H9WO8wKpAjoibRLyT2QTDI/YN24ujcli8INj9ilE6MeUU
5wVML+xFP7I3RjNQAV2jTMEDtd7dXKiA63w1DoL+7W2S1GssGhvLdLseSbD7t0Z8lsfGBFjniOKC
0vprnm4bIsdJkdCE2z3abUVqHrUbZUHAt+O5sd9Cy79VvVatu2ienN1CYkMXSAgGrObEmdL6aagi
Sy40cLCRr26cUpSPFyUX41t6XmBRYQmwREPRJAZcd4qMOooNW//PDG0aITpdJQ2Zdv2Gx50YjchE
ngN1meIe5V4+f77Cx8uGcwq+T7Wp0D0ImMO2BCdRxJP6a0LpuY2Itn+EYdqA3PguYdMbnMcRd6A7
Is5xdMM8OcB28YOiCUQiMHapG9VgIrEsj4okMipdFObzSe/IRzsEq8jK2VJSPjy6+zC4h5yEh6u/
1CUqdSYj3B1C2arcP5pDQdTV8MELhzETDAfTwawc1PqAYi4HGsI0HmG8NBnXfk3HzQ+GrQA7LbSh
IxAEMFH/L+xympIhQz+h+pOq5/w0//cf4wZY0MTFvXdg5FL9n0MxwLQY0I4NGPaeZst2FBl+XmlE
iWLsZoYIrFk+wg4qCAIFyP3DoVJR1LCLpDnri3t8x/wIQvUdNgQn218goqno7lZx3yRXaibL/ohu
NdpKcK594Y7J2ohbnCql4cG/80XUHWuGIY2YqYhjADYGJsgd3rp+vIdQR4Iy2FXvLolRp9b+qTGE
8LmLLGzs6CoSV+k3YlOTzuB00zVkjNae+jnRVxzaSV3Kc/NH1o5KNJuCc8X2r2jvJJKAOqTJFIsw
RASRwb9iq/ub/jW+KJsJQjZDzd9gf8l4KPSKjmwAATFYvCGNfm8fefUnCF4BWOo1EcWbLrZP9xAD
5LuOgjmenrQT20m1KvCl05IiQTocxSl8WdxcQgk+jAtk7R/w9O2JNZup3gHfedSyHnwSQkJqMtUL
o/CLu3pohSn84JzAmWhSACjrzIZqqdMP5IyeckziQTH/YuFSi6Ncrv8yWexYj04fVndKDzXeRiJ6
Y6iilRn2tIITSdUcLELsM7uaGBT0Mey8Jllr0Z8iqm49ORdYlSTAWJSChiPJQmcAVyK40+xON+p0
Q2P8WpMm2pfSiNHAttvl6FCOK2KSVOMymlswG4ywSZghzAw3mr/xs6DFI0O6qmyIj4ctFG/5fGS9
GeZw4QPVq6qLT9w9Cvjs61R0K//2IlNG435JtBvcbdmm8hT4RrA0lWargjU8kd8GLpJ9oX4Z4oSS
Bv4tN6XsOP1/0w4q5tE4Mebjd6UiTNm/IgZxnwj+moxmgUTOlFnlRn0BSHlShGZic7d5Z8yjSY7o
nz9YjqrBqktzPiVbFaEejdod69bVKc1wrJqf0oHcmtEhg4EeBV2meLoD20T/9w4ht5HDTox95H2A
KmkpF5Rb64vJySP4O8AaIZabBXgOUNv8lilaYqBNdlKg0rQnULMTJUIskcRM8Rw4KDGePbOXiERx
2F5PXT9keFRkgwCQoEu5BXM27Ekd4hl4dbHWhdB8nDFXrVzY9opplWsgmefIIt5lZh89EEH35Z/0
DDSm7bDLqX6s8TTItpsgvO/FFGXtZMJkcZLesMLK38tDfqbRk43wib7acdJYy+KIkQ+mYNOrsDS/
d0u9L8a4egq+KwU2wl6TCpXzEn8UzQNLoIN/Ulez/jvb5xKXH8i1OBLfiR3k4Z4UhkL6caEllsXS
kG22ODtFkwBWE/XZo074yPcR5TOjqO5lwTxqW4RBZeCp6O5FXzVL4FkiT6yHP2i7PJIR27gf+q3g
yfkqZjhf/Gu/pX01efaykGJtYcbQnSF8fdceTLhzp7UKGCQJ2WW0Jm58DhmO8Fbg7vocUvVyG8mO
2K6LrjO0P6RsFkPKKnU0LoSUhh/QkazAWlBpFPOCoF7LqmZ3iVHidDwer618TAJtvBlt0O5dV0da
vvYMqQO2vILeTeOxc3Vm9Xi9E7lBK3sB8Iu+LjcIa3UHy14EkGweHpzGCKZaUiSyHWqnn/KjFSv4
szGC8BhYrZXR6DtfU2yDroU1D9kh3qIDZ5GCfFjfRdNqbmlLwod2u4A5RKQFdn/0utVUYSDN+3SW
zJBvrxeMdCEheGGX+mNawazauMwqAXMDiYzdTADEkC3p+2bynqLxgAbGz1GTw0ubOUkEtCDWKdeS
X62JjsjPSYm428fBBR4lDt3dtifjjx7Gv4LAHp3zBx90ecv8YoJQiKZ76Yv9Mp9hxgejY+EUkudf
yTlN67qWOclIJNw5bScZExwB0idlW3AdOz7sAN+qSwyDmH67u0BjmTUrUxo/VL2CW9NweJPVL9G1
VrsphV+UukWaN5ViPJXGJMiJsu0b/SArjjeyv/6ZNqGmR0qLRP3hdkyMXSULXCkjOq4td8+ruqqu
0UgeOzZRFqU0oLMcuKwwHGW8/ZbqyqoZo0jhpoaO6GH8/JiLQMfx3nxEG0syTBSDI38Vj2/iC8So
U4z3D1Y8BRD8PEPz3JGjgijed8/a5VOoLePIpgjUxe9OFUM48863nJF0D8hqaCmNt6OufRiOFrzg
62de+/2kklLTUb3ODwRWcMZBjgXJb3Xwfu2Ofky4PBbQt7dNK5l6FXCskAqxqoYc9oj2J722xod+
WgfGCzyEbollI39CjSaAPRIiTmPUhChc+rxf8UWEc7EVdOXyHkZnYVjTuDIJ0emp1pKwM5cBrnmO
0lyihibdSpJZ4oKXKKNlG1EHlSylpPI9BFhikmYdA2b/SwojcZS3duvxiuDpn0Ya4idIhQRXKHAs
Qm26Wyv9MfqS2yAPSXCVpQnobYM8b1hoofaJhuY4bcOPRekbJEQAoxM7X7qDPzXJnIkx5Trj3ZeZ
K8r0g+2G050IDy7pTOpUC+ox//Cy+pvQDUla9BROecyJQE5nt4omTB3hAYjemSEkxQ9jlND0nzC5
2Tb38uh4AqQj9fLCD8FdtkMTN0IJyVLkuY9KkrR/YDTFvUxUAglnt7qcfWWd2AmyD6WcneJ8rd2h
KyjZ/XDZ9/cVhxkLduII1Vcy9c3ppVOw2n4p7pGOK5xyJmt8UncuvS8Gnq9E+mquAOavUtuJIPbb
l/0TOdWbjeFSfVRiqnCtG0Omg7i8mRB/Hghrphmm9x+BBd7jfXElz9sMSlmZFdFmnr8CVhHavA49
CT9szQBZzODMNRaZf5z16jlX8WBGQZjfTyzpVfQU4hjz+gRzCFolxBpb1wUtRqkSElIHUN4KvNes
164md6dDuMMkhcqMP4pIag8PM98WvEdPxch/NyJ8jzI0xDv4+GWmCvm7oZodM6Onivoo8ZxDPEEr
4P/l+8qelL3YyON3rVY16Yi+RdAVn6YYLiVUkN1fscM2JSqzO5qaEfllFHbjdfYUUA/zbHD6impD
tKoD8Axj48JDyewwGaBo1XLtUEDbRU6jgqU5uXq05qUv+NnAKX2a/R9EcfjNuzCF7EkbcDwsXO02
EsicwTHKm5yka+892v1/UhmC36zMInkFZXK6td5uNSzP9ipTt5pYTvfNWV68EqBmd0YJsdyunYkk
WgzbIgez4hdzpMRAF8nuGHqWGWFBdkb+bXYmER0MKBNir21pv4KY5kUsUtTqbqXckKN0obNKjqTm
UC42PgiQdaL7AasxIhVtOJRSggjy1cYK66tes5URflq0njmwUCWLfqMyhr+mt36wSDfJOaV0ViNC
8p3surLOjzyS4NfimoHP/GnWEOV6RlVUaid/GsdbRAClg94RaSSsQTMI7liyYA0637Tj/gaq74Ik
nsvfBNY03zOzuSPFGtlLT7DOAU5FH51d1jyV3UR3LIrzQMft1G+E9rWKF7qI/eWBq0cPdRjy0QaE
64IU5WDJ4/rEOZmz/evVvVpOJ6PuxjO/02OWqhlqE+ej74aiH+TkXytgFnTdPOahjf33AyraNdt0
aGKteFwhxGDKBJI9Hjs2WKUal7DjCUBYCO4aHS5ka/phb+LboCR02v404l97XCtkep5KqcuFoGCx
9mvLf94FkVCQL8KLTPMFzt3xRtv642f35+2ZhxP6pvzkLnPvqHmv5u/aMeHjEtvrvwi/Vviwq16I
BElOcu+gu9WrLQ+zrKg9Lsglvh2qmd1TFCobym1/dmDUW5NPZ+eYjPDxQfhNaXV+VSnQ1OL9iDMQ
n5Dcw4pHJj/gLepJ4Y0HRBIiR4XD3PR1kwjH1z2JR5Gcnt6WpTGWnU3SMvzPmfsOJIuSNSitCfN5
vtv+Szd26GXgtLDMXu090eAy5bSjKV8xOrWp7c91jNzDNo8veRvwr0wFW/egAYtkx2Z5+PELcGrP
vJhqQ9ZhnRQQ3pMSiMkNccwFbmGggmSnsnvuW58YxBdUVXKxI9DAyOdj7ADIPcr8pGvziZ4UVBky
reMX7CQseemVkoY/2di1CU3RB1KxTHSdfrz3+B1q/b0OOOF5CoAAgLYyhkwGI2AL+QK2Gfoxm7Ze
5QB5ezLb7douSK8snNmAGm0gb5fvct2AlvvoRfqKSR61ewsI+qEuRw17BXTpgUFaroIYx01C6i3G
v74zmQczC3BXZXHSI2OGlpLGcUGlbXxQxhRpd9JtOFQHCvP3vewdgz3hJJkWQDEmshRNuPHvIPq7
9ucFhFAQ2xHi6IrmF9plWAlvHDixOeN0yXxyGgQQm0zPtZr9x7kadkAc30q9Ps2F/dMfunxMg7uP
BhzlIjIagXeBe6gHjUkTeo1oFd9WtwHWg0JYgCSDIXiluT7x138Z+Q34oLHZRfsJVRCX9aJ4jZNu
xYMeSO48mxCc6qWKIOyTt9u9eRc7dfmdVUP5lB5+hvkjzPjeJ1Yn2R1UANDElv9/DdVEW3nQyYMc
/zgHOEOWDu6J107hQBTMxnU/UQa2/2vr19DhzAhHOie+vtK8tWOvOxq9NwXCOum1IA+1iOKEdsAR
J4khPyINZfzAgTmSwUC/FjUuHCCO83KYQqCujNJ9nNS00XlFxxYzUGZr0t9uCtQcgItHg5e/TNsW
2ROS9m74L9DPxOdZlMkcNVs2jdzoSjcSNWYqMc/w5cdied87TAZLaR5Hj/Yl8k98PXV4KyZeisU9
aCGwRJS1UTD6VeGmk9wCgtVrRdHzaq/VSaOZcbjH8hwWXwwWdA/x0KSrWrHthTLz49F/shoMXJbC
gI/r7m2YFCGo/Nd/NCcYWTRRiNgNE+5l8RT4xT8su2zxcTdIu9sO9zsW9+lhEamVgF3SL8DlY/oD
5oCynEmPIrgnTcQICEHAuqaRX/nJDA4QIWkNM/kdrWeZqqus/Skcgxueg88L2ON2OBV4daaKJ15W
x3q7uhbiCp25G2wuU0bF4nqxHhrycRCZNotfTW5dq7kN5rzHCtdVbApZnpi31nV1piG4Fo/x1Mt7
kc3FjcqKnrrGb5TUSvOGcVkBrGSQuLKmNkm3L7nHob1PMUpzfnxeIND1uweYulF0W/+N4WkGCYwd
A9vlRg3boRiqay9dmlEaxEfD6TLm63+ybBTG3/VshBLb0eMdci89X1ojbfPrQs5BAsTDbXJdSXV/
5f2qLgIV9fpSeXe2dlDM84s8rNP/PFo00CZdtZZbRYjRcOJTWFSRY427sIz1TBeHEEzbcltFyud2
nFbOWL0k3gkZNzAa7CnLvFPIoCydB1oBMKr37JJZRwa0iOm/EQ5g9VisBBMj2f5tvl50TlvqfcA7
Sc/YOL0dK3J4tfyH8NErrY5OVSqpbT2yngGmeRG6q0jBHo9D0qwommhm2V+xTNw2/c5aEb+7wK3R
Hv6U0C0r4VIfR6cuMy5ZsIulHuUgPbENmlvpeaK88M+HPvpQM1whARCmvg/SNY5IGnbc9Pi4z8XZ
Pcdh++amNp0oqgcLwyhrwRuxP+U+k3qCDm1OZVj6/pBreqZVLpPuUyDrcK+mTs2WeZmpE+8e2Fqq
ZyygOIyqwyLShQ8ZFgj72meOi0+eVvtluYuaPANxggizB6gHHDKCq6GIdLOW2JjO4JCyQKr0peV/
ZHjgvDgOSH+GTyqzlU1wJeYPalERiPxAtvUnzLHVnIKy3RZqaQi+uUG1AMMU18u5ok1RnlvJ1YcC
b/Vswhu2rNeqebBDQIz88praYDIDsBL/42JOzbSJaXoG56WWPDZ9bfCWj6cLkvX0DNy2NB+9IR0h
roIy1Up4h6V9lne6OTuxZN/NdIgVfvuVhsap23JZewol0eJs0cGLA3lSVvVl4R5nWxw//Pt2E4aL
xULrHvG7Vn3wW232XUvZjrYP8OSkRsQjIH1tIYXz65Cpy1wNQq17+2ec2qzhdh5T4o+VLE5tDlVa
ap+enFXAyWo4ZTY30P80ZVTSSICcyuekCXHrRM/gjknIlS32MHU3OdK7mbUpOc3+nu4dz12HNICV
qxHc96F4LVPWPQXf4eJJOJGUuSpHpkFNhqX2Ei/wAxFIL4JR4ut38NwxZi8vgKrch7vi9qhkmxu7
ULmQ08UDP/iRz9PHZo/X44KWBVzvfWmvcJAua5sFa6yXnkSiNej5ayrT5vitvCggkxbag0n5T1bl
59q3mdiSQKoeLIol1KXDDWJyxXKN3U6W4ygzVnG2WasDCOHmHD1awgyGbHKHZPdP3ER3LAw2CR1o
A1xOdONNV9CikDgcPS4JfCWeInq+nInip02et3f8rB2TChvB/EyFWTUGBfoxSRTu6SfyTgR8Ol4R
WkdvVLY5aY0Ld8pOy3Z7pJ2PN47HdYLyHBz76BBGPXUvOA5oCJzRi30mfyPgTiKLqfs1AS6b5AWr
TSXU2SiApoMVzrgtW0c99ySI8zg30johVsrlZbu3/4nWKDu3pOUp0xZ3QA1rDPLTetHlec2GtLeq
aP8462AvucTAYH+Tf6A03lofML5w7f+cKqzbktMKzujfTqMLsyr90fY6Yo42b088to77ejxp3Blo
N84Gce86g2vAJJigteEoV+sDxn8zB1cpU+5b3IU4ZX5tp3U9YrrjmoqbDobi3lSnn3Np00zJ6d0S
4WdNX42VrBsmskJpy35QEQuueeDPTxQPEpPMOae4waubUIRjd0Kd73J+R37/pcGZr+RuXMQ8Y/2J
pe5wpKyXZC5HYe6qIWAyuu7zR1M5j5LNz8vhzczDuKSucmW09bd3HU+bhYcS5l0Aa2x62a8wmFon
Rk8cqRDuW8fGwI7xgd8j8cK//CSZjGQCWOBP0daMYbrIvxsewtL8eCG+/lloqCGjjh32nff1erFF
+LnfqDKC9vhAmvvEanomby3lS63WTaAxo8dmlzoPPAmHAIQRdTgcztPB0+RwPVSdUJEka3PShT16
8pTOYf6FgSTQH3cjOti043BnuRlZalg2UJBfgoMwkc+Qu88UYChpGlqfNgUHxW+grKXrst5uXapf
7a20VDZV/GPb7PmrOyv/X9JVRdSqv01yg/uDeCwWP0XhZouJGPPz5BnuBjD2OwckRdzT7I6EHD9V
Jz5kCPDQH3OPaJ6mCJUGHSegcWgj2TIBqYHaIzirVcUTVJw62peiuhEVyyNXsATvg27Cn8TF6GKd
FL7J2lMIDgjKWJam++7es3PcAz1PjXzBlmnpqXr8vRS3aTyVqaKavlPVVNXPjNXEXL0Q/MHObeGx
2bTHalEoSP1O+jmw66P3kldA5bMaZBrK5ei58wIlxjCxgGH9vtcQKj40dgLVpIN+5dkt18lk0qMX
NetdhIZ74HZPbX2MkhDwEg5+TuXMbx5Wfqb4saeJLixCLxxGTtiUMQvLRMj7yed8MefhXn29y1pY
bUq+G9ZWbULIwL0/wDms0EDyn0T/SVZ/cGJxVOmLpTLmNvVxxnrTSqn968wFPoeMhuXcMMl9Chr6
J1tLFanqGfpOaAcf+hivo8t4j8pb9aqF/Db4a1zmFJJnGOljIyWjSjDPxG4QFE8eVbA7BM245e4u
YPwp5ccQ1z+YD0FsTIQkYKgcFokvq5PUYoNXPb9y4iSkwanV993pY9vee6xLmYTtAq+cWfEJIyan
N9kn/k1RZijgCNyP7xy7bcauw+AXdMXptroEE89yVHF9xNePtCJvHRmC9btWthLZ3wtJEScqI0B8
ZrozP37jbHQ7gcZwRcUe3AicfB8+0No+mA/yVnWv3rZVI6U0lperdKSRe21sqmONJ1s2lMmRBztt
SRS44GYaWk4V5vl9prlexgfmoICuwRfk5w9kmLBFcMW3EwAVHVFwTIv1CpTsyShY2BfIIJZyY6ty
S40RWMa/8XijhJ4ObFby0e9eWct/kjIlJe6S7C1mbuvvTR9DczSsSAjWB+AJk+Donl9RoQOV5Ksg
QWUAzZjC7gHF/JupzBXU9w6WsemBCg1UQvy9pCISHmSdM6a8fezczJknNkhKA9mEKmpkDhyGhTL0
Uz15NcGhRiN7ZSRqOrf+bKYZ6aYDSP2TjwDMtnhELkbnjqi8cB5LvKIogqF+cD9HrMpshkGu64c0
leSTSqCd90NlNEq/t1b/jgjrqefR3syGJOd2x4l3AvWu++yc+YjjXVBMV1nLZJLuX7b0O3jxH7+A
WiLm2PrrlluYruYpSaje/QoiI682iyJcOT0344yVU1a8t0Ldrdp7eylhMcHeMCjk6KicXWqtS6pt
2eUJee1ANVF0peJ/RjzQICB0NP/B5n5WiYqluJFLFXBjDiTZBgWGSmUwd4yZ/GMtgSX4hFq8Po9y
k0gXziTY6alvdlNx7nBLnqbAsIz33Gr1xID71gvDZuHfDWatfhuEPjQhpPaVQJ5/ugp6m4rMToNI
WWWMFwKVP4I5fkv+0TB052Fbl9T9fyTLknlSNzICm6wCis8ON3iwiiA/qDtPT+d1h9eKX2wzCEPF
UWd6zZOyS1Go2ff1+Oz/oIL0ddJqmgbQAGdpC9ku1606DvG0ETzJkePXft8K717kGwE0sOSP1fMF
go4Mu++/34nLHJSgaZPwsuODHPpvOOREiTSo2PIA0iJJkpu8wWRL/1q4/V1EZvHXZloYA/+W01yS
QPd+Op0Z3gAlyPKjGL+mRXFM1q8/SJdJHKvt2qWpI1jH/Xm0AElw14LXtXfxsk1s2TcE2iFT5Odp
1GPmMS2EjwEEuHk2qZqUXJMCw1RNOINswkYE41bKgL/DVE2YrN4+AcQv+QONngHOY0/RMKwz7N8/
IDdokrfTA4K7nkueR3+2He6mla+2W21VXRgS60eb+peoaMZmQLPggn/Cwkfyn8b9Re/negWMC0R0
sYpJ25uaHz1P+Q4qA2Y7T1161KY48Q+1hzve4A7Im8aSQYjEvZGhAS0StKpADU0RGljxiMYdYmFn
2ErMXYQ8zJo1+5+hBnXce78y5wMJxetsB7XwRSYvnN+w0RrE4dWc0Lc5O9FomrujhB5LpImsLZyS
Lgr7qZdgOKgZCOBo+wrcgVArys63K1u2wxgPaXmW7JluOlh9a082CXkyhqq/d3EA6qirdVfiLomq
Eb72pJRtIl381cKXIYPv3em5uR9Rq0T6FEsQrkZfq+41QV3Uff9USBk7Vf9roBYOleO8A0kKCy4t
LYmo9RobRj6aiWskxZ2tl8SGumJaAIkVLQX7hetQxtqPTG+5X0Nf+Ln2eN2aP6Q3UjiLQJL1hZG5
8a9x2AoMA6Q0FUFz3UG5taAo+tCyNtWey68gyAObcZh/yPLlcqMbkHq/w74zKVmf8Ba0mxDstZIJ
MocVdHLf4vtXnVR/TU2eCmO7fZ50iD9DJybJ6+F2CEE7EG4k+Hncu2lNPJyNmZfE5Bs4Jv5QlTmt
pz331ByqmwXwiEDk0cTbAQd94WbMKToJ3LL07J2gmwk1+zYGd8bOteXVoRRv/HE+aQAyOsbFuwoV
K4MN/iKFadY14v0uG5pWRX25mRQcRrUY+O79/sFpRO4I7MjJGrSsf+gxxeIJLIK87Q+Pn0WY0Ulk
8AfGBRFtSHGxl2EhSoYU+UC0f9rQPAgMnkWNICMAH9EA7GKtzL8mdGdDJhLYCFQHLGsf7OyAzktW
YwOWKS/fOhzrGaB4zD2C05gZ01knd+mTEUieDgSD0AD+rCt61IYAt9hPyJSC/GXsPzRs3y7G5vOZ
2S08fZPdx9XcCfXBydiVp2X02q2/3lRzfuE9nh3vM9XmDg7PDoobchrd+Ry0ejV1/qQQlFeicX2F
16RpzflHABqsIm1tlcp+mHZJqirZsJId6r2VnEJ4jY9wbocVxQfK9zej9efTEuSr1PhzNgO2q8Ek
MTISGzuebIkMtllvvjs4uE/yaAPuKNnqyGQOfj574tomlSchU0zIrQDa+HOhLF4dNgoh0Ym5H4hC
MexhdtXYO3V+N6uTWbnFHdwONKmO6zxqQhruxiadePSRCl248Ys28hwjy5lQAcIcjR43HUNZHalS
zVlXHxWymydSPZ9QRDIbT2FVn3iInaJ/oupNz168Ueff273jNfeThn0FppqPFl1vrTII8snII4bi
+IfJ9WaqXyP4YX1AxAm0Z2u8Dd2YImBIa3RN9siNOlOuFUeDsoOXJtzbUkBTPbTKSRn+iPpjWmuj
QTJ2t9ODjGVC0CNs1k4GsHPASHVeZBDO79QF9GD1a6HjZUt9kf8g4OdqLYZvyNah9+IsfuO8dkb+
fJL3mXDq3yHuv0o9Mtg1V/HV1OTUWmIseAR84Rfccd9uBjc2v+KioBuax92LRpQNUyg3avkwR1qf
lhlgX1chLL/jzLj6utAl5LaP2pJxe+s2Ld/l/03kktwwjLAU5qsrp4E9u1LbbzTkkSmOgPjfeOcK
XckTCt1MIJE0WBMa+QgI8OPiFQNhKyQ65CWi4h/GIf22H+c3IKqaLNLjwxACuL/TLxYNJNVOLtTC
QnVcUPm1VOulyOEV3ifldd8LxDp/1Cf0Q0xkd2dtDHIq+zMeJL9MG29U9KOqwtvtnalyjrTcO2qe
eDIz1fNmAT3mAsFVUFH/HMkT2YCFZ+ucoeAUe0aRHZ5tNonI1iSNyVnSPXUVwMLDY9E19/Qcf5xP
n3Lorh/uZBYxlIKpvCfs118sKkHVu2C6izdWAQhV+Uf8+ivoqqxg4cct6Op/mYSKrDb/6hQjXb8P
WbUA43p0EiGhla1MgYDJaSCe3UJmTKRtP3aRzZ/l/jxQtFSik/ugW63Q7RGrLULPiluBFvX1q5ud
hwSbOKebAUTOW1NCkMIuPgzZGCr/rJHa4uQiXlLK4tEAMt0ojLbn/pb76f7dmtIbpaj0lEVKj5CS
RUXpdq73FiupzcCWhTznrZMsvY7ZEpZzI6n27hroM/D55Cgo2lAQMOf0qLOA8omOdWNBRFk4TKpz
Kcdf0dypj0kMr31uVsi1PsdoLee4YL9liEcUMtBL0cPatpMr43NT/DQqn4XSUN22LhE0+TItLBHP
UEw9oXwGyXsHtD1oV+M9c5Wbz0pNxPBrasfpf8Vc9gQSXEBLboPXeuHupDzq5KsSrFjjAeGpp2Qw
gTQVHCIvaSchJKy+DRpxfhFa9apiVl1+mNUBTl0tcQ1aivg08Ot1NTS4tJejca3OzxD6EmtSZ4K+
0/tN+UhZa4ZL3IddkYFma43pjGMXVWohGqOM6BkPu+xiYri5hBBI844JK+ZeNXfQZ8brQM74mJt/
4aoIB6MZzmpZrf3DZDhhujDsF0WWmDb0QwDLEfe9ThpXk0AyXZNU0bNLNmhrbPnsY9+Cvu2oYUi+
W69oaGaXQZNWrZVB/DFIAF/OurFCbOdSFXT7u7GTBlLQrcuKutokpYaMtUNl+sUvLTGp2VXiF9TW
uSN33e+YWVtCal6Yb61Pvv2hAdvJ3Kc99I3IU4m1HG8a8jyQUgkAhlEbNYl1K8Z3+FEUwBlqgK5N
3uVfXMDs7sprcgrUrLeEHUt5dEHf9GHBuh3BwJdxFgP42bs/zG4/Sb9MUdK+Hx8Vx3HyYbxCpfxy
+0PNBn7pkLDClvJ8qbOb2Czy1GKQhf8JUm61l08WqUuD+1019MFIK1c94isQToCE4KGfo7Ow4BId
0Fj4fk7dBOdT6WO1gPBcOB1ZGqUN4lPi+eN8fnsfWS5nFLOUbnAGo25u78ikJo0H2Q1kerP88nGP
ubeILiWU9kpqltzdIJuw20YNLNqB/b2mGEEdOYQizbOpTH1Qme7cQ7STbeq6dC7WsEdLtLvYaQ4t
TNZgGwlU5r/4Bt+9Rlf/awwSArb7GPZ47aml1Qqa4XyaqGjIJEtS+pWwtPy/LaxJaCWDGpzON/b9
sfM4kBsp3J0Xwo76vWRlZ3YOp+lA4KVwz52WCD4C/K7BQSEmD9qVw8FwpKgBOhEg49piTUE6BB09
53kkiJ12C6GkfXupODaHnp13FZqkYcwTYs0hR/oX+HUl2jhIs9LQ+y1Y6ZoFvlME8qgpVLD1I6eA
FgfHI2tItZK3giX4iiPTSv1khsEcA7YaPV93rLMIFnXtMLLkV4q00JqnCsxMxgAO69uLp8QljhaL
PWbh4IEYU7lVaSU6G2PEUyhYBsmCs03HVz3I89wvDrB0B/GdThyI7kU8XXe74rkN/eCoLyRVSgyt
ux4YU7yFjvv1IOVYXSZtv+prvROhBvtRPYKbPea6oKC9q5biLlUUpeE07OjzonrpzMmn3NFtqQFs
wCOhbecT38JUyumvHWYjzU18Gk+Zj8PU6T27XY4dZCtrHXJNceapf74+iCvQzTV+JPVGW34hra80
u3gabClQBQTsoloVvkJ7YeEBged3cdw9JX4H0V/S7g0GE366u13hv7LqpEv1vZZ7K8ZzKwJ+onZd
qGzX8Mzte6K8w7AQ7R0bRfP2Nczzo5sh5BGtWLkXwaQBwu1idVm3jG4rziHovmVyi7r43GyqZ+79
xnM7ZAmUUggGr03+yZDmXSek1BB2m2Olt2rrG1p+IgqUKny9VvA5maeRtk9Igqlm403WPRjDxjle
Dkj+EHqyuUP8TuP9MkxuCeqTeA9cenc8hVsXPFDpUmAnBcXGoYBVjhUB4HFQZvOrKKNp0q3AJYXr
hyv6oFJSLcnAngNLl1RN48XDQSVciM4m4m0JxVaKoRq+U4UUTcDKJ1hm8794MTd+qdiCxmyTErnM
4q6v9JMz6s8pzhdcbD3q1liZdwWqEH3OhU7cB2fNPMgG+0Jg5dt5St/15VmVDoiVNQgGmLIZbPHC
tIZ7b5AaDYZprSDw4jkRZnNiPXZ10vrp1ppUCvkL9SC5QOGWiws3Dz8nVc7m18WWzYXmjSo8RypK
cxCrhxRYtEOBQpiznWgo3JHhdRRC7vfc2cqT6BSaHjLYHbhxQaa8+IKU4WcgbRXCy5YC/yUzCi0r
M0vOZjT4XMBO/YcbNi9KsjQhP6HgmPU0gY3pHvFVNpXt5vnpBz9hmwV4LUx0JNJuzyDW+g661pLM
gRVfQ3j9ElZ1pRJR80CgnrYkls435c4JseFu3PTAVgGmEnlLWHrp6WpBqO/29zfAgBXvIsDBZ1pR
T9pMJnD63ar78CCqYgxiYe6aL9M42MZcwGJl5kGQzyMNf3NQjVTroMSWevVfRrxVukdJL1N0/SR5
P9jwARXvhq4S/Dhp00+bGOHVYSwn4v330Pwq1RAeSaraFNg7NgKhrvei0Y1HFJ+Z7HcSLiC0WMjI
2OX55NIWOCYP9DO0UXd6NjXcSRzHcd3P6W2A2ZNUTsll81I3YtKUvrRrxKIDFg10SXD1OJ7c+cG3
8BIFOfYma2WG3FtKVXVDA6m1EI5508lNcCSCC4Th8zyFMssBErdoqYsrI+jWWd+Ibq5c/vESAd8s
1MLOE86Q/QCSMnVMi9vT7RPRQV9K7S0yfqlsssdbC06ZuMdGzB3nzBqa3pt4YMFainKHDNB2NRpZ
HoRFAYH+qDAk8nfvA0z7OTED6842jPG3larCPWn3MElDXPvrqdCONyy3WmxNWXLN+G/Uxwqrs9+b
TF/X4XBDOsIWe+9deZ9DH5kQ1dQEthKSjvUfYelq41CfuAu8B1mdha/pvGVWbMzWHKIaCzXaGmcc
VYn8B9vT4KngsZftcRrLG3faRR0uQObbSe31jFrpFnMTwWbRXa7Y1MB4NbqwufrO9n08fHX8EMT/
pLlUMsMkWaRPwJ7xEtg2WMrE3/BCBK0QTpjrRUOJj+AqxWtzsKkdX2LqyNFd8q3YtfZ4NemL4mXz
cVcVDbOhZN6SoNs1YIpQEqQEeJSbvVH84EEZgJRgkPtZa5t2QQFxrTSNbdxkNhnPTcBvYPkZ6+zU
UIBuAIDDIfLKtG51n2jiaLbDPoYy1ahqSrQiCYIbxjgpwsDyeDCV9NQePDJOCCkMiJJPv8eND26y
YojJgmJJpacDEflj+CmAHg64GmJ3FL2AOjmsQjIEepexkEn1FDfN1zDXHdOy9O36raMlREWdRD/+
3u6yyHTqjcb3GNZKqHZ/e4J2erN7r65khptEW6L9WYtEraAHzE4wIB5i4FC3yL/xhFpNbtX8AEEX
7FWPJ1QTYAB7KPiaGdEYDezMRBjq/yRMxPENkaODGt2oEJhLYY90lTDPtdAiq9hh5G17JgKwsGj7
e2pYEGGGHQ5w3YsAhEpP3D2FRL2N7/IXlrOBhL9TD2uoKEqD6JCCWMxZUCo0BFFQKcc2fuITTb7U
/rxp8OByZ3/orzBuIjwdn1uMfuVSoSsQWdsVihbmvsGt4Vz1hat+KicJsZgxA12y+xfuChfGp3HQ
DYGZV6xtqy8ZIYR8rCvifxXUZI0rfmT6kNA9bHXMK2AUMOv8KFYLqEaoilWGzFKF07YsExtKiy5M
OrSrfwvMDbdsP53Ps3o70Q2UT665tAqM/VAJl5V9mwrtyDPkfNSnvsTX7GdikNEg9CDsWLpuUIIs
7U++f+3lYsEEHkvLfSNCdxOFn4oA+uEDgsMTn945IAnUwIjnBHg7ijSp1+PFXSKi5Lrelv74CpRt
cCQW9UBIpYlodz8AYGFwLnh1dZysM6fvpEnl0BUr15L48AOFrx6dYXtWc+A5my/nqLBOqqLctoOh
zhBDG5FzHgNQUEnCEHcQHZEsLGm/tuntU9zCFv1ny9gkuA870DhBPkVhnM7otYRBnzLcazM1FmwH
3P2OeYO3Jq7vTS8BeA1IlthCig3jj5x0MZHYPbnJQm6eikKfx7giP6Isbhq7wfXN0S67r4aVTqeQ
8P2GHDqxmRZ+2v+QEbh8H8isgPPJPX4H3L/yPbB+KgIMZw93qxti+4mBS2r7jpJrrRIO+1+/qfYM
rMzzCVe+J5xo6bKJkfzzJEef0LTYOcRv8Ed8e0CBTyYArY5l63OVWEXgt4cZdSsIdhhOM1Ubk1OK
8gAF0D5tIQfczWkvkU3LjUX3NWr0EQWCs0DZbDoM/8RMzu77Vv7QNijObB2pdrgzrJrNMET+KlCT
nFsYKz8rSRot1dqY7fd+cZrfB8AM9i6p/cAtfmXVmDmMLtmRJSCunlMI+j/DwGD2Q5n9nfkXhbmT
em/yXwvxgVgnoyaI/z6oMHx9xgpy13xm3UONMhlGapHJeJruPOHX7Iyni7qLijJXDTxZVlEC5Oqy
f2PyhbJ2l1DTRGha1+gjUZxbuTwt2HUqiSn9MrWXdHZg61Y+Cj0LNk9CNFfp90J50zq2fsCRqNsP
Z/nOHFfPjBHHsBgkGV3NoUvKaB8JxICaeIuoFiFRzngAFWTyh1RPddaiTBxjyXL9KHPX1NKIXYig
x4Ox77Wd9ggWkmQYxQAXfzlthd4GRKxQFj71XBRX1Rr5ptV6YFlIiIaISOiXj9+CUebJtG78PnUv
8hKIXedyAgV/LwsMRmmSAKRsfLvoXq39UQ+A9lV8r6suBjHGDw6VZ9kdygimJJBWtpAQ3JM4tt/V
4lFbAz98GcBjswpdLUHhVmdIDGFJrWJt8NSLoW2YUtpX/g800IFzT2nDXBmNCw4ybVKQQYTZcHpR
qub3vyCoUY37ttdcpGc21DZQE8d6jmx6WIkbkRUtPIBhITG5p76p1SOTgIdliMdVdXu8n3B+toEz
KLvEHU9WRWrsoGtOVA2X7pD2VzIz33aRoSHhMy/fFlHkoQ9DhJp43ZWym4ReGU5DJurZoLlbXhSW
EijzQtLcXbfHAUTNzB+max7r6C3Cu0Ht+frwQAjqqaQGdKeQ07qhDOi+ILtmpVA0tuSUZRjvcog7
2i3pwtiIROcpQMkR1/IUhMNG5B1f43RiiT1kgoO1I05ik76oCHrf99yR7sN0krvUiyRzKYp1iwy0
ThFdaLMDt5Mj+x2NZ5u+8r0nJfmxDeAL+zyNDuu8hSoaFKFLjeUC+AHryNb7JkqPfwm/wj688uKl
6P9FGRw65cdWBQ6TS4a4fPjqfBfEqUeGVtileegVHK1F7QVit661dSiGxUKgh5b4mRl9qvE9Rlfb
/c9W6QL1RQn6qnbR1jYbDc1cyVyphmANCsC/cxeCR6rgBc3zFTuTnjnSttKzsduK2GJBkHxG4pMU
ryT8BSL36zfg0P5/fhpcpKB+8SLDgeZeJKBh+0+mT6966tfZpvXmGpAde/ObRNUS37lCUFpYEkuK
9ur8vu62jLlsMSX1enP+QMoCtqvuGGiUTEc0xTXLHL0KudfMO56pMdr+gXV06PZZN1qpugH61jbX
QMWZVr5gVb8hhedafb6FuNp4FgXfEUZjBQhONyewwcPif3sDOrAYYf1bPaVvoLU1XwDPnhlxZ6+K
C9lgNo6Get//z5TVnsSo1FWtBK5IqZPxli43GLs9L9LG2PvVBgEqOk+0p+Zj0dHToJMfe/w7w1xQ
vxM9bhPGLnMQRRMOlF+iakUcWNtfAzaSm2okJRr4nGTCgtzMM7NjJp1Ub0KpJ5f02ascYK0mNAif
2rmj/HnRBYID90q+3IQI35g3taydlZn/3nKL94+l7N06fV2ajJ/5zPjtFOHws7S+fhqnBVgZXVzd
QIiX4YtBylW9tfZZrGWmrpfil/YBItexj5dRfosz6/3El939xQ7rFm5g9kDwT5/oJ48Nw1Tcaq2U
qJ9P2JxjeTo5iiTsF0oVWmCKmd8NrhvYIEhlZd1mdyGGQoKK+fBFEWJAsHomi7gCfRL6tpVGbEO7
Poksel1+G7ZxXG1MwqPHnvX4Qe1+O6ruUQ+8d+saxeOsy0dGJA3AdTtp7JMZPnHQYqM9qGpQzfFV
UYW71dMcyoPa28b+H32utJr4Pzgxi8viYrOW/sesOQWSZ8bjomJ2tOwbc2pneMIm+BXiu5dnm4wp
+YcVGT+gxMY0PN06/gJ0VohTo9NMn0i5kILc9pfSDaXKOMuaFST5Jk18UOsse3WrdfeTEq5LwUK3
bMdZghVZDBqq6mKcClJSRLJTwQO0jxw5vhJy3keAr3/OuA3bfQ4aSGt5q5kL5ffHC13xE++0n6Ul
3bljYKbwtzruAS7Z+u0P8SXD422tSdeiNMyuMtMwsPmOkAA6dYkDeC4F95UjAGJFD+lQfqCCecTC
4p/T38VBz1IohiYypWzlsw+mth63iXWbIOvxeP3eWR85F/nI57uTwQCj7LXjMHd6k/kAqsX8NeiK
yZGAFk/oWCstZxojOYpVLse3Dy5ZE+LnQI760P4P9H/l6TfZY5iUt0M/wNFtbu63NzJg+h+RVoae
7QwKj/odlF7z72ThDdLuQehc8FCFULZQ59Fs7uny+hJhfRIW1+NfMGbhW8hgzAEZy4d7gxioQ2oG
V4m3VPJvmsOd/IlQv3LWBEBMi9AZm8ehTv3zs5vvA/VPQt5sYa4gnoGWGLd8pigAPwXY6dOW7S1+
D4q11qCfoLEe1ESBi9MmkqdzbatcHeRDzvjnER0fYQgL2xROJvkY4X3f6ffSgSuLJdlB2tMkGV3x
V+TTMBRlArbl0irEObsHn/ETFf7v+grx04jcUgUzY3GG7GWWdqQIk2ZPDI0UFprwSW5n5PAkFlZl
7G36KoAySpWJNWnvWq771vbO4jWigH0H++0q+kGLO69HoYQ3SjRolXW4Uw+MjS57lNQ6/I/20gYv
ytufaGFyTJvKHILjF1dy0Qki/gS39hWfz4vYWhl0H5wnLY5XEhH+e1d6R+0v2Kfq6qgMxtuaPioz
/5eRWuZI3uLMEiODmxa3q1O/IdRtRfP3WmYKCSrkOq440ySIS2CLILVzDyLRuJMfazxOaA7RPQXw
NEWtLiwy1rmLBCrMCTGYhbcJ6POgNma7DQAvy8YQtxQ+oRXBz75A/t02u9DEzAfK4wIZB4F1Lb8L
1aZNUTgmi3Z1RbYX+V6B1fBYhBYt20IagJzrCtdfDsBbh0kIUIfP+5R0QpokUry+JKyeM7TXJiAO
Z6bloYUxfl3yqrFtyu6NfCW4kGyby+5X9CIRBagnZrRC2RqRcGOs+csXi1KSAouWQqXsY4Nz1n12
ywXDxVunDnzOUb3GUTKkZxcOciK85CZqBwmC8iZ8Xd+aXfCiZNlNlgi3yQpNfvuaWI/PcSm9Hnh+
r2/kujwaSc2QGxP9HDHA0zCMire3MkUqSnCYkWZUZCetg8S8gxhjp1VFeIZ6ULyRbfdI7pMVdFel
2cugRg875ZwXPOq8ZSyUMBLb4US1mdrVLsbleCUpHhwPYGX+PpwVMtzxXBxWlpQJAh4ilJ1UaBe1
OvM88FNHJOGw1z781nhTFHwe1m58O6Clfm3GNGv0yTOnzwUhtOfBtLgAYm0L6RTvhQw+PgSSC/aW
LvGrcwLg76Uw4N/9XCvouEGXG+5z7imENwFYiBHcvs0SUnMem6WtKkImLAbuy4AW7UUVKevG1Ley
mSVpjRddwuJhIW5HkVx3bur2S/sgDvyIOevKFkV6mEufwDHkvoFrSZqLWerNgyDgRTGsRAQ2pv57
UG65RIEJD8+8BQtS4sruHnXXNSjxFwa59SNH+sQgdtwjLpQZC47f/wTKvJSLy6EFerXdcbsv19vD
2NDBbGKgff9fmHQyui0E8MdIOj/jP48UhpFrlL+k/3/Tzj6NMeKmEY2INyNGTTgrEC87KQ7dnMmG
mNR2iSauePvvUkzTPSLRYJ3KCjnE1VqV6Xx80NAYjleq/eD7Jmk6GU95PdBhusv4rIpwokHzeRXd
ezRhDuSHL4SU+AMKvX+C414QX3z4sauPRUIde/3YxIqRYJt5yAjz0md96wkzkyPQYClcjDC8tDQS
6cY+mdtH3afLWfkNm8mzpYbAZ0XjwNmTrpKmpsjVFLyQdt2y6F2mCyrGYePsFSoPI7UDMAZ6yGhg
5GIFMyC8+rkyuGPo8Z5Zmc61iuaeFlBg/uH2qHFoEFq1v6yMfiASEFN+jWS3VJDLoBNScOx6vFAb
U/zs8pkw2oPxe2q4zstP51oHa2hYMjcb0NjvGTDyWWD0/qJPv/hPjzsz76u4HcsYGE9EqlwrONo7
R70iRQFTcPgpk+8t8uJKddMm6RGpFUNiJ2rt9z5Huh+iV4HyhHNxtT54k7hRHGmju13lAoDnLC3f
xKpTVKMjolPpy1XnxWG2d505ZGpTcrLo9YxcoFtkvrZxqZeWD8nA2K+m2L9fQua+umIRrnSkEY99
tDDhip1/riLqN9AsSUS51yrPksqhd7f+9zo9p4l6q2OZLVwFsp3SUVko1mrLOO+oB3iit/fm87Uc
1+HTOzyy7XS/otURseCI4hozcRKylmOIU/AXOb8UmrNi1MSLe6e2hDUeCBhlmPgPd6rZcx9IxTpN
d2aAnS6rbmvudTmsCcqEgX25W6u/cna9bPanJqaiC0NspHXzFbNt5M2+SbXcjARDUT+I1nPXqFc4
eaFKhJOKLbLBElhU56NBTxTET9VfjG9qreFjUD0Mnfr7ULmhG6pkrMgPkQZG8QmN+iT7Uy8EK2Um
bUdxqpT6EeazvNtoMOh63QkyeDtd0tUWZMdl/X8U6JKh+ttlcYlGcsYxmnDki03QAmM0FpiCVU3u
yeq6htvr+ERC9do1g7QiYP5OQWdKIR6eCNAfL4l9wjdzpLiEaJ5Je/bC5Jr6Ey7pVXWHeyNksUm2
ozKvWDK2qjal0B6Hy6TOos3/1WaLQxHEe76US02Rt5Z4QHqp0AZsmSMJrahHbiwAIv+7OTE/8rrC
dPQrdHQj1wb9f+tkoPmMSnXztfS+K+CJNJZT2v6kr/f5w2iNa158E9LXdPCHxIaw61PQNss2Vsc6
PofZ+oykh+1MMcc3qXUmF9FtsTfhLYH2o9hdK5gVKnejF692HLEoAm1iMgEO42kfzPkNzRVdS1ko
oxqYWZpRRAcR6wtJzRFEu+yR24n7vTOARZVc7b/Y/2nAO4UuGr31ku9XrjZvUi9SM1AYvKiUFxtV
zGiNMbLypyZCE81HBuUa+GsQuPzUqZmmmlPHtvW76BdjDvE1jV475L+Y+r6QRy0RvO5qo9z4wENy
ibGgRdh6R6sU22C/EAhCUqBS7odJnxuyTWniXWv0bTonRnXwPpEq6zECsC17CF6OyvaNhrn/+JFp
WDa9Zhk2F/sa5pSj2t1ccqXH5UH5ShkkpLZkccM09MGsSDvghRnIRGuoYvMkZHby141pEvoX6lal
1GML+GMl66qBp4Hp8SOl8A3zwhOWqB0xlTfN8HqFfEkuo9mDCrAdijvFzEjrtc1AH7quUioNblCM
p8ZMKqI1Wo08A7kleEigXir0sJePcL/DkLHu/IKDKcg8zLsFg/0IzTUigFH1UdPVoe1WHVwTusvX
QTzVxsFxrXzwZIWpUy7Xh7mdgBauIt1nNpqKsPau577KA8P+E/h+w4XX8mpFm/nPBfU2YgR43Iqo
QyQNgrX+XsLohfTHS75AT99FY5yKVUutDag41e+a93w7Aj/nznRtbqrltbGHQn+y10QCNZ9+Ox+k
cBomxhOLnU8ivZg52O7s23xj7DVXy7Ft0yUekOp0vDomdcT2yzni2L3baVxe3h7ADmPx9BiropyP
GPs+1e/OVvibCtWBRLFEF0g/n35CQpRhsoJBh3dqpPMc9Z8hWH6oLEZdjmbdPGHxH3fBadeRUuHw
RSC1xXL2sX2EWEgyBhYQHzy3+VPE0pOV5L2No8hl+6A9aFioZ/9BvHhi3IsfeCKDRRMzrJgp0gTD
q86i1sC6v0SblrDV8+n+DasQ9WBGifYR3xHN/N5naSXR5d8awciE1Dxd7EydMIsnxFWuS1/OeObU
bJafXbRwoLEzuDvsvNprESHA4r3TMu9ZKn4TvqkZOnWIr3D2rL9fo0hXBGhQqq3aDlMs1iu64YvB
RZtguhtduPcGG/HyubVLnXI4KaWht3gtQgS+ch+MBuW7AGNoPuLkBr6x27Kpba4C4W/G7/ZR3c5R
7Jv4zyWL9IOK+CR1JNVY0gIAG8SuciH7KPNadsiI9PLAuOASOEOTxqlbHu77pI4BkP5NB809yncU
MRIvpaJ6r7vpfMkci7M6nd0d+vnI1c/FmjZUQG2r6WtM0iwzpdQuhahBnd/dfNROFEwlfv8gZcPo
8UblKantmoNHIH2UV7jk3NhwCPP7eOWV8tEPVqDUe5+w61bE9trHacZZsI460i7ZYEhJgUQKO3sI
KNnnr3uY3vRmaBiHvcsnDQRN9QRJf8chu3RcMqWxHytSESPgvzVNtWrQ5MWfYBIVyLtq1qqPWjzD
8YDL2mb8DgcfG0mrmWsIZx1hfbe+4/l6aX+l7nMpJeaR9C5CHRsnx07//nl3K5ohOX8NJtvCUQHh
Xa/RWTzkV95I3NUKJv8AK1cwqWJC32QLooiPP2IZteH5Iz/vANOtd1yz2Ot/bfp/C1yiKxNtXm/H
vYe7rz/xAvOGIHuDvwqE4BCmHqGWhqlNho+lgBM1b7hrhn3kIio773HoQqJVa11yIxkIrGFyeFtE
0XTEkV9+GDgGQ/j877Mpe8xKd3rXJbsjIRev+H5P8u/It41ZhDTdmJ4UmPFpy2Ct7jMn4f6Hy0F+
YJfabPotnm6YPXcRYf8Jb/xbDF7m5G67xZfI+3Og63qufbwMbyjJHc+dXg18oF2Ng4RRLlzrsPte
lHHfnjYWmSnizOlpBo2x9uM4KyDiRb6LNfWDC2S1vG79ICFQqEU/EOR0LnvelSmhHesCr8h4cCBg
ULaoiZmrtqK25H6KJ1OILksYnjQYqtI6PNgAUnPFC4s3QUs66PNs52RnDe+b+fN6ikjfGcUosaKc
ZJ5/fzBRzjTq27jxnNh5g6e6vd7VPVIUftPMd4GIUkY7jU3Vs7PvGGF+Frgo7MXg5zcl3UxCAP36
Kxw4+S4JoYxkMNEvsMVE53j3F72syUj5kRoLTL5rC5OeTmaVNdpT3SezNpxldCCqyJ38md4aWtEO
iiTld/Jx28o9ldcl8HgdIxfdc6Pi/0mfoGntxHXcOdfQL7g40wIUH1YFSMNWHisGhdcLzMuoKSAd
3kzIO/h+B+6LhhzLZmFbs3R1hly8lwjDxB+l/B14VsEZXY+ZmPaeum2+MreOHd5/hZOAKRQDiwfA
IlQ8cm692zAz8cdMdgg6kSoLzscL3/mnKAgPT/CNtxm3IKfmkUSa6ceIJfBLeefsvVZXvf+QlGVV
csjhSOuM+H9nHn33EiYV9SwGK9tGmA/42pG2ATpugHQB4Dbn+DpFlLUNvqjTnX3bzKvGHSVDlnM+
hisQoa1J7+d7Xcwp5lvwgmKxIFZT0bDebxi8bNkaK+dE+QcH4cIE5oO/hbofqb4CEWdyiTOSRVY1
7vrh7gLqvwzvkXwbAUb1p13UF+Y+cs4QF7XtBb7C+eheL3eX6z9SsNp3bUV2h6gCiHqX9/x6ux6h
lDzbcf3pHgDtj8yM6VHxqJmg18QvN3VWruQhgYchkzbFzEmuJx+Osk/9MJdSVXsg87Si9hkKIvkR
Ri/VbJtnKCjjoTyoMnl9X5HsLVkLBI6asEbI4MrAYwe7SLkO41fZxRLODHrussj3HkEJXY0MGTSY
GjMuhgxe8usRDEGJCjjIhAmvP3k5GMs/keXItjVZlFH4aBlT8N2bjN6BHFKhqUmF8bi6WbXZlJgh
hnvzCpj0kLZd0jq9WdOHqoBN2zzToDrcGM3IlpJR+FjDIKBkK6m/+JBTqhur1sHlYhq3rxrDEOWg
vEsZNOljObchPGm6Pmv0FMp6DBnvrCRkUFAGHqqxoBU+DxiN2vz26eFHNZD6H0u53caXs16t8xbL
ayOvF01NPwzY1zKLIbXtuEzY6yecJ7n4G/gaXCANX/bqoAWDl9gTFJLDE9XR55mqylv9IfkmLE6D
78OS7dU9nRDGXBwosG9agiShLVfhlVOcOBtm50ny8nB9OmvGi2s1iWloFaR1es3e+Jws0ZLOcY/Y
LDknPck3DkEIs0vFte26L5/jbeDcbHkbyxnul+pK65appeadLIQo6rW0XKBcC/v9k23ZYykaP42D
g0r3eXVj2UxcX3+4pPsv3biMRtvDv7RrUowNrl4jC+l4LBCSuYU6vN0aAMCkF5oI4KPLLujeKruq
Ag0fUCxml51u6B79CyIgZ8oZsC/z9h3GTLTIl9qad2HEld+i011lFrFmz87FKnCp7VcdS/6FNsc4
plBfHE7fIWnhrw03t4XkZ50EIe3XGxI5mktvckHLutr/bhYB1eMKjtrZs2WobmFKSxXvsb+pFMcn
jRH/Ui1I5RLsqeEXV0wlyQrH427sr3e2qrR3z6J1UWeWfI3s8d/hP9ieBpZ5SfrWjIjKhSkjYYXo
C5d5DfSHPRML2fFvZSVzGQK+zL8LSqq88U0Vuw81cPdKCqwcUz63e09SEPaUlyhLWlSoDgxEeoEv
p6fN/JdnbR+GSOa3hN4gXk/Qz8fJZV+RnRn5LCFQxxYT8Ivovmi5X7b4asr1NV6J3zXmXPDZqaKE
wYW8GpXbdmSUDnuIto2CuhLU4CeZiEeUuZ5Pfa6IylyQSg9BV1p7e7ye1zLWTzmlsFfy3JhMft5O
bSdnSoV32ff1kS9595ObNT/vAuV6jkA83c+S1PzxTPEYzVOuaCJBpxdnECD+SD5Dk4xEq2Qrdg8A
S9kiziX+a5SfqC4pwemqyNnVx4fVs5F4NLiI/uvoeq/C7wL6A/Lq0lrjOtD+0GuDM0Ez9uL6N2CI
KuslHhfQR0HQYlPT6BjFRADWsvtbUJY6dNhyVpkrZTpwkUAKPJtBjrxGcXWN6mGhAoxbg3Th2UJc
dY9PyMB8dVUa/KgqOH92xMqtiUviZo6zHNmLNcAh0X4o578kMgGr+E0Bz33Z7bV7FSAtPLwbpT19
hkyLbTIBIusCfcLeuXPxdfPXO7bHu6p11mS8mlPGH8FsVPeR5LaAUEsf12N+fFCiYreUwxzwSs0P
2x8XqnLHjMvEy1iIZ34BTdrylwZN3DsdIAt4OAR8ywPDRD1ntMdB+LHwi1TYaJ4PgffcclGuP79N
lcbqHP1rf0n3FwqIFTYBX5EvJt0uPibRz2TcBsHqD6T7rrQc0iPwHuqq8Lmklo7AZAN5NfZ2AUfa
Qo/YOtvqNEwSOFUW+5OQu9e3yeGUpZwWQrTElU5cP6dCq7S1VDDoYgAAXzTayrYX7oYwYnmILBjH
HlaSksP7tsqG4xfURFc+NbUlkDblrUoqj44Nd6PrwXcR2Da3eCHWTzQAlcgymwMAZPMQwQFq+dHy
D756zBoJYUyftzcGdZ34dxztqNl7vgxjylf048+GUaR3M4Zroz/emvvF2aKczqGcoAnAK7/5gmnm
KdiF7cUeBWcHV6g9WCCjyDddiW+usJMi0cr9WIAKsTTvbKyQSRBgmPCE24cwxEO6IEhrtiU/1+1K
SkgXsYa8ZpnfHZ5YX9f3hFjRj+Q3v6vxWNlOlnkhh7ufJhwsJS3MvTkAgOhhCq6mXX/YAD6urV+C
h2mfI0bFVemaf3Gy0mWb2nBlbYU0uFTadOWIgZUIcbxmhGYxDVMZJIZTs0i6oqlCNSKv1EbvIpm/
MH9Fe2XH9kI27q7aW/TVjVQqB0/N78M25OZDO1JjHODN/GagscfvlY9XPbGfPQyNpHKigSf8yw6c
5S1RbvOG22+IiwJblh8YuZV+eYRxGbCQ1IT848Dfff2InnPn3rITmFU7HB8jyHWuq4UVeSGrp0RQ
ehNoKDhTUaGune/KJm58m+BhX6fkYKoAVv2jR0R+6sXdv7ZYFVDp1PGxjCtUihKl3+XSFUj3NMnZ
dYADbIkisyfLmn74OYZa06JR1/KegdI8BhZPQASE7UoP/47Jd37FO/iOPJymGKqae635HKRC5PB5
LvIfI41IvYBjYSfqp8bcIgM/eERKwa4asOl2iYkYWwti7J6QXdBNirAvr1fBaCija4c/Fa5rcaml
LuRBLysjvWZfJfSwGNqoNMeqzdf+6Y88z54uIOU8djayN9hIFraMpIYhhqxuDAjlnwsYupQsv7pk
s188cLvs6v0I855JIn03UGtvzWEcxTLIan5AyommUkzyUTWcyUAe06lUiaGPwmnvZDiANwfqocPr
hXFSVkIPaW2D1Px7mAGaqRkrE26Nxe1eRpmJYmzo9T+3adNGC0AYjiCFUYMEHjuFMLJn0FIMGdww
od0KqJXChO8+8PlQzAGUfBFpvcORkhP9mcodeVlzhjfn3hV7d4VZHSuy25qwWqppFFF4PuM5LLg2
pjuV3Furf2FjGDsPdQyU1limxD9cdfv9loeq1kSnMcrT9NnlEQQaKKceXYjEDREEwalXR+64UicI
o/vF+1XiZ0a65QiwBrz7kvtiUAesC4GutBuUNFajEaBuap87Qov0NfzrZcTRYmisU8ez2jPD5nYH
jmCbQHcgpQOdH4Tv9PguuMA4T77R8IwgVg9MoXDi+4fz22nvVP9ZhLGvjKrUnTneV2+p1d5Oua3H
MQ0QLuTe6T69ZGlahjcahkTerQVJ/JbXyhwEfA/w3rcX1bcxo6N5Xns3UH8isebkdxCJs5oqP2Ph
6X5RXkT8hkVntoTpaGr7YyZBkcfdDKyl1RShy2XXP6E+T8agMy745hb279O9iyv7BoxSlYQTVFID
0HYTXJRnVu7MKeGqKOWep84aa/lvEUNxuwHfoyD7vVG19rYZ3ash7XQQX56F3LehTVVgtSl/bhb1
M8135NJDVOeQxAqI6jkPQ8U6wMuZJxBz+Bv2eQ/TcGFLJU4mhZ4thLR9dZ8LDGCeO7p21Lnje4Vg
VFUKD4gimJauUPYsdysSobHcsjhoaDyIa/rI2aFw2EGaTcbonTRP2tG71lkAYwbSyzr6UIYEUxL1
omymyvuZU5g9xZHYDi3BhCHy1tiiCusrQ9ekJad7fBIEI9AzdyQZDalCwDYSeNf4yB0BzMQuOW8c
T+K02/uBd+snJI6NNwkctz7ZbkpER93CTGC8y8XeIeGMbLkEwHAqnne8DZfHjPp0XEH/1hXVlHyV
Re5VvBAmbeyqGEfRANL090AUOchu09wSgWvx83aLjWVdjpGgjn6AZ9c+tYufmroHfcRezv3wEBKC
Y9yDkzQuTY1osLOH1yTjcDTWUFFTUcMIGLPLh4p+5nYgt2zERST9PjEVyFKhyu1usIklUkvK1Ktl
QQIPok1IsfMjaCDZsbmrM2tRjT3NRP1bVLKZ6JUQg4xr6OotJleCQH/7NcHSm00WRveTnpXbtgRO
2YfwOGRKBLCmkRtM7Pd/n+jpZu7psuKNm09Qogw0sczQ2Ele6k5aqHZq2WAdrjwClDFqtgfjhfpc
mi2aWqWn2A/bsw07vrfFsbWBLXXb58a044bnnkITldqd3BrLI9jD6dDmcIP8vTS93rL6VyAkuo1i
akHrlLxxWb4NGTWwRUZ2xXOn9jLlrJG0wW9F1m+rRD/RwvWASn3YdwnbAxiEgFmuuNYBUqiOOsgN
h2v45gIi4N3jorJZsH4pmaup3cXAV5gMRey3Ud8rMr+1RJBAyPjRtUOvbvXvUdpscDws0+yGl5JW
GEwAz42WSdaxFQcacattHcHXJvrA9aGZ63k+h1IsQaO1z2ONXZyfQay/fClVpKQ2gmlXltB7D/Nj
gMvknYJhD+onIyN3ZE0h/pJR5BgogwIziVHsWVHs9WBGQltMn3+WXVFenW9ciUV4uqUASb9Z1zKM
WoyN6wPLbJJQ4auq+szELbkOsdM8CaNxxUZL6r7sPylcxXu94DuYNarvw5PRu9l7ZNOgozleq7Pu
aFQwJNw7OcW3NGbbfJ7eIC1wkynUC0gXFF+M/eck6TM+N07KmzOZkjG5cehFhq0I6jHFz2uggkzC
87OSFsURN7Js56C/AQbtWrJTM4ItZD12kUIquZYq0PrjHDng76a0AG6mHzfc3Mptmp7AuFM7pnDU
8PoAmg7k0kYM/zDFLudUrlpllbHDN/7vqa8nuXyERj4LhclfPPFrh8iMoaNtzXWtU8KttNLdlJj4
5EpH4fmKO4gA4RNzxOJX/MapRHgJqrN12KvvEhLJaIdX6evng6bqUt+JFtbFeKXDrW+vsVamhST3
0mbmF7ZMCoVF/BAYv8h4gjekKf4a1kI/GbatOOQzjHv5MOxSR6ye1s+pFjDUowE9iqncVwP42aKs
pvgCIUGBaviWYHGysFmkvoBWxxNbdM62PscQlLIJWD1VuuIg3YfQDk4+pmIU+CdpiIFdI6R3kiHz
8MW+ns3ldVx1C1yE8OBTcKDybc21W6fp7HyMKDWmMo0VFERgcPk1GLVJuhS2TjS8QWGRtnJjDNVU
AJ/7b9byXmX4KnNXAtUcgwr7OpCfXULa9MfcWDyxopMI0eKjmc2Ddi9Qyb71FAZrqQbcp6u8+amT
X+vZh7S6pjjVsgHNB+Q6hBj63XqtnFPnnjNCYu2kcWX6U++r09tqNDc3OBE6drn0kPjMhZY61jHe
B2hGKT0t/xGSta5NSCBUpe75I+bCFpTJR4XqhN2LvSedkwym9U063VSk9BTgU+UvhqlUjEjY4K7O
iqLh61MdzkkqgTJyqkchN/RNX/3z8WtQ+DsxSUPT//sfASofOcJi6GmbqQt6E31LTrNDsdpzxvAo
0i5D3HX/gu6ji9lev+/2YNgkaiIrs0oqYTeMyr9za0YEtE/BQYnwmC6fnzCAKpWqlJzb9EJDV8RL
bFknqu7Y2UIvIHvpW/6Zm1TA0QqhDlfMdYIqA5LpiTL8ae/MXBeMLlmZOtko7L0aIvZmldL3GdjG
AjmfjP4CtPC3DyB98X2D9DwgpnAcUVBn7jdqFVKvSaWE4F6eT6e5q/zg/n/jU3GSHym3iyTz/88W
U7mw90huh6MfVFFYWKLEf23KHHv0EIkDIjg1LxI4Z288W6Ku1ptgCENANNahGWtdkmUHVzA575jt
ENHbX/tF95f3y9HI8wj7tVMjKR4pUsHbyIBudOXrtTy5rWRIok3j3Z5jG1Kx5XCkNaxuw8bjIO6r
qpFiECuK4AB9KgGwSymowa5AIjpNDHIiCEYBhGNB7jjl/xrMyd4xa6orM1j5BrHBVAEts7IqKi+G
gdO2c+kJakaCvF1K4SkvluBGt0TwquL5BjYxM1xoIgEtPCfD08bQ1wvjK3AtudYVRqaVWOT/bS+0
DlGcXqCvEpYxvtQky7xNf0y0RIiqP58jgYsDqMn5fhKkr2ytuuhln9jg/nQ2YHIVhCzf9+Jr/QVa
BaKnfLQPhxZAlbs/KzGKB8L+2M767PqpysD6unZ8M/1zihukQ8p4TOzWQJGA+YAeYeORi6TpD/Cy
9JvNdYUrOPUoFFuRItPq6xdLQAdaHYvjv3koM2DJ52IzBWpywML98ju3LL1XGqIksK2hSCdYJnZ0
yeIyLIuUwSTBzhjBuK25wv3uEJkP9Fdu87gmRakC2bes5CMoALreIMaid/qj2Oa8QZA4/l23hfnX
AB6VEzadViaKJFT2kReFyVpr/n693RwGbPmw9huN2Ce7N43XTWvdSa57Z2MwsvcA2czN40pO95K/
TiwuTbhF8xF/c8Dbp9zsVd48kTJ06ejbdLYtD0K2MP48YjE1LIbzaMISMl2qWCdDv05accu3AHMa
52+4ZHS+SHxE3Ofgj4fmGHwDNdpuwhRUrBe+QgI/zmOMJk7IlfceE8O07tszc9MOhMSt4+ILoODE
wSitsedWllZ1+5wm+HgIx1npR5u5vAb7pgs11JLZDK8B6rkdLviBVGXkgWzynxytvsYqBBAQ5c7M
/8SvzFmb5gUykp83FUUAuERoBQwveFPTllsdQMe0BIiVL7YOAcwJQK/LB/c3AYmP1rAr1fhXJZ9e
pxQbWdz/I4RD1StiH0/iHAaEPomcHLbpjhE8bbTMi4UT0KQXM/neReS8812eOr+juBMyacJ5WQt/
EUBGbeOGSum0BUlZY3BNu1Ol6QB+85CVQn4JeJcoNv6u4YErvbZHdnzB5R6jyQP/raN/XjtePc9+
qOsE2n2Gt59kOptUJq+G5s46qWWY+SJM2bWoCLupvaLVT2n+zc7tmGOv17wOHKxaHwtUzHI+cHxd
k0llFP3TNz/PeiMPliAtT4KU+oxSPJ+WfvSWtXdP/ykY+W2KiolcA+TKmV3vpVxCqyC8tmtHSXzo
MoiHBdlVsceWN1F4jEsFo3MmGTybkukPMe0NJ9mBXzWvVOYHvd7I2CnhNFAsJq9sRLMJO9oHtAkG
iH7IEtK5nL3fZNM7tNg8mKPETk0aFd9bVYCNK+CF7qUfNzpYrY+pIa2M32Zd63ApMVTQ48VxWpYj
tXMf9jremYOMVxwy1u2Rae1aCqooxNWJ7UFkpkbV5Vo42dKj/E/2codcOtrE4yojlm7oOWa+tp9n
QSKgkaMDw8OHiJ2f2Jim0SVNVqjZVpfweTovthB3E5Hl6CQfwokuFvuSY4lnUGyKiX/iDAOij9GP
qhDIbyr61DRMmgf7rm5uZ27+9zolRl/Lk5cPhlcqoHdJC308atsQQy+v2CAzaR4PqC8GaupvRpx5
xJYTQYwHnW9FAl2L+6XZ2Dmt4Q6NPefvah0zOaISICja/RU62/jxW2UeIaTzpyhLsQor0DpvwpFy
QP89NfTkRKErFy77votMYgbsiiDeoYlI3PjlO9FcxIpIpuaPaXINQ8NOsXVgCexs9f2tsMBhjPG8
oRtdEgHGMjgBS6K8QbBYOK+gkpfk36Fghwc/HgZkweDGN4LRfDEfhnk02j0lGEVN+AZTuxsWYb+9
noJKofyyvXkP/ti37gR0JNTqCzEgdLQcm5mmiRu/5Khp0gAI0YgkzkdXZja6PqZQ77jNZF7aq94H
rNoj6ngcw2Znsu1df0cwrB+pAkh+CIuyL5IFDmH+czMr/Ly6fOLerj7HeDiMgVvWHOx0xbUeyzUm
HHTmqSBC7f1/xW/y/v8u+enXAaGEmPDt1hkIhfr7wIeyygADAyzCXx3yq5mjnN93X6cAq1VSRpSX
nOdrTm/ZKQisXRZrc8pDVN1JwtqY9sXV2/2+k+UvUaQ5qgx+FFCwyIXcopRkaNTaW/46AIvijZ6o
Rk+VqQfHyEzjXUx+JpcF5BxDPPQoHAMKV/9Mp8OctE2jGVHYql4nR0edaYvzxeW+CcCzgKaObamv
YJUA6gjE9ske5URxuNUtgibXBt9F7BDNCbDCnn5+h7Q9e75SbcBxXkqo3U6hl2rRpVfbIwjDHRu/
dzV3aj9p20JW2x/HkLDOSZe48OQlJlAf6JM+x8eRPuwWvSpvUO8oBN236kucTppAEnB5N1tTkKK7
W+ptJzzJ7bBLfg+VClVelSNle5xpfwIj8zrVTn1fdvpWZH6vW14GKa0MLq01pSa5aFNn1lKsCX2y
jwqlPXjc+pVeSGa/3sqcY+bA/EnV4ueIpiQ73PIXlQjry0bm0F5K/wgb0+i61WIuuBrX7TuRggc4
bGQJosTug38Dp+Al+6pAqks1ecqrgBGe92EeVfjrNLCjIEZBEBrLaJyjz7XqsUcdXScBMl0AYBh/
eNzvitZ3gCUedE3NYV7+y6v3RjrwcTzulFXbBDO96eX4An565+hHUAv2MfMnV1ghM4lKIXdm/zpc
eOAOUAO3S4TfNthg5JKUTmer4FrRK4ZayIuUafd++xK0UNbmOsuw998vl06D+p/1JjddLl/9a13s
eyn36E4xoQPVWiLyQBwXAJjDBPV2AItWRo4uYHH9kLCdXNeKJ3QZxTzgyBgdjpHXUR2Lir2NJf7C
+ivIaFLQqMf1ChFANoSqbEkTzkKzrxG9GKchkXnCbZyhJDwgc3PYaevCwCn1gsjIkBrbBMgihBRo
f5HQueU2fChOB+JDLSZLHpMk1hSWf7P6jCbA/twRm5PWlpjkH4tg+5SXeA0CK/ef6Ut22a1G7EvC
6IphkUHeMdpJKx/Mq4VkMJbbHV6G7IGXdRxR/Tq5qXInfGI5cMrErh9NVB30LKcxSKhX8QDcvZuW
IjAYNButjE4Vi6/vghTq24/C/oV/8skrDsqwI651fhqu3LPpDkwiyUEEJ3/83AajOaKrpCcCbbG3
MfFaX2rv4ZyOaa1XaBGCVSLkoMsmJwr75bYdeM9UdYWq9uUS85Rhw0MrJkuczZnOIGh8znbjUwa4
1xIaAriLC+A5GT14KdJ5gjbw5pYs7dGuiOtzeZflvnn0PK76dZN0qhC1G4Z1AHe+dcamqLsaAIs+
iRDSDKRZxCr9qxP0uzVPxLi4DPuKpNJ4A4hlM6klFgpmCGoqN4uiIOfO7uI6uR6QVXo4cDf0NyAO
G+IxUjRkbaF8rTARs8wxzkwnoVKErsauQTBHplkxg/4eBNfrh9WHcjXyX62Kah/tkK7H4Y7mIwvR
i15i2OCpbTzb83k04W1nQjB4bxSPWkwsY9FRAYx3/ESM5h7CDdvqzUkMLNdqrl1hMp5IO+A4ABG3
4nZZxLy/F3Ui2dgzknKNa7cFS8CILD3R/Dt5LiQxZs/gNGBda6Z7vX9ysKYJNMyTEmghs0u3F1rn
qYCo4DCP+HxRqWNoPqZudhlnJ7A9pfs6t2AVLYUhauwWQUhCKRcozJ/LseC63LwkYM8I7Y/Nd5Jy
fEkwXC0MGNBPp1VCsI3vG/TfvcyyfBScEicZqkmrAmrV4oUvOcYaSaJdJHSy6a7IlaYjgs6y0j55
Fa0c4GKyiUP9IJKL0ZrxxtMb8ThvvEq1fdR7z4CaHpAkfx2A8jA0N5Esf1V8d7t/Pz5wrD9ocDJb
xuECjmBjyeci7biHp0TqExALrXA+2znAmrzIgiOA6lu3B/Yb5c6QV8Q0Ch9zAEtdHEXMSEbanfXW
NqiBdTXqcrDCUPCrh+72bE70uJzDJjZp/94YV9/a5k/WUOZpvYOkqw9fjUFZQKaixnSHnbfrkfXk
9mxHIdkAQKLWs/o1lmwAYTN7Z1vaMVvJVLPTy350ZCFw2cmQ3BbieHwtpz7WFHdHDIG2KG5R99E7
Kc0j1+0DFYYHkEoRD2iHasWji7ly9FOzn+TOegnwD8nOiibAr4eKFjDwgjNFeRVO/oItEqDTrGGv
FDKPmOoQXM7TOQ3tQBr0PWnugmNZyz7JvyFWw4/vhXt3L3JPJQiqfPDWn6dJjb1LFthU0wZlhlRT
8mvq7oHBIVPP0oiNC8Qlbwo0t6Vp1QM+tDToYlDUTU8PAA7EmmSqHQwpwOvwEVNVdoV/tkK3U2w0
PCW7wJOZ1wFyn8YBUdhE23YHe1E3700+f7RkQyz11/6hdQvriEjAVeLBskhgvlYSOCfWfusX2P69
Zt5tZJ1lD8fAXDKIoKnUwwe858TVcWbuzodT5hsvf8Nu5/H91zGFvrtp+xFAxyiHROpkvYoOz797
JxZ6VvBGXaq4OYztqBpJc1P+IuayycwLfn1uKrLfZbVvExeYVO0I0eAXL1J+z+nLVOHINsODm+Ih
+C+MAAIUCgQowJu4DYEyyXhOWxwSMjH9LAXFL3v0tqPYgofN4gywnE2wKfZla+h46EJssDK6GCqm
NiSzMdrbab2bjOoIc1ClLU0AtoluiuLfaE4UqZPrxpHA/hghB9uro4ySg9/WIYKEDk844lsl534A
W3TnwJ2UhrNBLiF4PoFWuNx07sd2VY4TLHk/w6aXw475uQ6JlLBARjrDisz6cM0ziAIRne0GEDi9
2d1fj5TFVa2+MEX7OMN71Pg8jXxyTlw6oX5bxsC1/PxI+E0mhIaJnAe8luvlK1qxysoQjqk7DMgS
DpCu40Zb+DfyubyA+jgpmXpvkYxDCNeqPLgWusUyJL9Xl/cHUBFAgc8ieAwEFUzR79AJcCW0WG3Q
fk1a4tHywNWph7WDVqKP2f1AiiKCQXv3ol02/c82LiQNbcfgsxgZXg6eFWymoZhc4dtz2HwLa208
B0WQHzZlks+iIrBOSkELpUeEzo0N/h4r12yMn4PEDnu6TEKBwmspwMYfFP71estqsJTlxWOhauq+
uUoqxFbWmSgmhq9xFW34NMde7IfvrKYZpdDugB8qRBnTCG2tcIRQF10ovAWZKLbFp9drspsbyAzk
95l6wrYSnW47lqmCQp18MignVVPukS6OAdDiZC2IoAhz/PqpbY6E5D1pDIBI5TOu0/iGXNsnuO6G
23lmScjLZBuGCgnDswDSDwuI/MGkRx0mpZ3lQs0cyPd8pJBGjEEwn9KuRkdejZsYrDcyPgGqRI15
j0Qbe9fM10fXg2Q84ylj/jouxesyoa6A5Q6+FCezkZOnfqgpmR33749IxkV1ZBgbM24numXRb3KC
sjzk3C6/qmpF9YFN46jjZK3NqHqcRpR3ucxBgurfKKkCsXqGeei9ZjhrF6I5ZxI4O00YGKWNdTB2
y2V6r7aApOU0fgbTrZ6tbEv/dbclpdlGdDpf/PzQDNhRLVLOVwuzB3dDB36t9iGHK+xgCDrdoR+7
MsLc6ocY4ZuX61FVLN70dU28HYrrHzcVGoeVAZ9/dSieI0da16Ils7v0RgittRWmZT1B7TIs5x1j
5oOTOR7flJ/iKaUxVh8SXZcmm8LXCLu7H1fuscdXBwWF1aZ5Gi8EQBr276SN9Nkg141mc8ysoMTC
/gP7CB54oprdBTzuWrER5K3q6qTvbJH6NqdgwOxRNAxC8W3FwbbcUU5v0GApPe79udo2iubzvt9u
eP4DUWkAi2Tn9PYQNgbhZ24ebSs0G25HaAabZClawHXS9gkjhmNvs+zUAtjUPD+UqHOYEOnG/jZH
kDLnt3M2U+eCScxwNd2xmsoWudWocJsHuMhTMn1rLG7bQznW3UJXcImT/R+42YNfk0bTwDUahWDB
DcEq9L2NTrjGgpiZiCDpwRK85bj+qq9HE5r6UZeklhKlnYld3mFuXbOcrp+dHnfiRbOIfagR/tVX
ywzF+PLrUxwXqXpwoxnHb6L8KHbqQWYCt87t61UJJChA73ImyukyReVzob+7XnItlD13uts1PH2g
sOdfYRRn3fCRfeC1inLTEp0H/Fv1dhtoP4x+YQFLiVsjdR3f0h7qWVhSk++Wy2xHqN3WXEHTYgXz
am/s8+mrkREKS3aqZvMB6757L1sKlub1ozjmqK6w671ExkfYfOffB858SNPGPAtimehWarL7HCUo
caTOKeK7hfOBcOn3pUMCUb1s3pp/Ip7aTJUvME5AA3IyjQHs2GJedfQVL1M1KSaC10b5k+l+LX9V
BiOUNiTOJQjvfVd1wwjd6B1eXOy+lgJWQL4olIcxUFsguP56YTpm00VqjtVs/CFp02im/tTkHqgs
JULday3oDMViyqwLiK2oE4PSnsynKMVUJ94/rpSJgyjwBF+4kpMPb6qnvJLWeTocV/u+jQbqKhuR
2xKswObVmNWyyTazRlrCCQH5G3IUjfYoC3joOqcTe6zjuze31SM3sf2JOJSVJuODyLKO66fqAeOx
fQTs22/ewKP+s0Nw+xnyBE+3FPfJYpGveXp5rCuVO3x8vy/fT0GJaGQV3ci0B+NcQLbrMieOa7jd
Ixsqyc7FyoTWiVYAwLr+Bc6MGL1G4de104knjRGaih4CGIeNVGPszcX2cJyQCwXTLmuBcov+zSAN
126UxyM5MIWjuyXG6BjUvRwdE1QRYonYTuoeiUEN1HUaVXzn0R50lXltj3sGzGoppdT3MG9zYvi7
c30CtOLWRxK0ALb3Sgn4cBKm3USuaJ1ND3lkipAjUUizb+ozdZIfq3AYmLgCOdm0QsKMiJqWvjSi
XPesDR6FnQ7z8kr2SUI1PVYltOEf/DIwmZFOnwVdul6qGvvAft8XqmpNiTN9Sd92Sxl/ltWZgLiH
zo7p+Nkhp+qqSKtcgboHpVwTbT+nFrF2RboiraxRjQX4TfWhBZkahVf4YwGMNsd3+G6W0wuQg0tC
WvSrYVb8p+BUyh0Gb4+/BEWZm0x3arIRc3r9RBcOxPbGGErRTj685MCbT4+8qVheBwfrnlNBwL7Q
2tFMkSIX66OXq80WB+Fpn15tfufFKmc0kGSpqQ0+2bEPgFGN6vbjDKJ7FPlfbyVmtKIXUD5cYh+s
4VfbZrveNviSdjxsVm4Elhs4yZZcCY2EEQPO4rk9yqeMDeRK1kPaWkD14O9T5CRsJmjIWPIovXz5
nFMjSwCMJi6/MbdtamOX6+xJ8KhWm9KPIDrobXEV+tZlquU5UD7eIoJ1EkF0Z0yCpit40lkV1YHm
eeA1FL46vSOdhx5ycfMMFLadaSXwXF+eyZEQh5yAK+/DtP0+jo0nRT1KQMzTFPd1cxFEmWhFz659
HYDJlhJ0yG9Jkeh2a04Pd2UaANwfEti3SoKLvwJoEk5srvZ7KyiWyjCqKiFkfw2F3+md5/pu+Dff
DjDKERr7JKme1whaiohYp/yI4hckWJTIy4qtt9RLR4ajwrX+FEmtos34j1xjjUOTlo1t/cixyyDr
LdJGJBsKPqgJnJ65gqGXQqafxHIGhTR9pp0wziNowhEDp6NvpsL4RX3ycdnoh8bY6XIXi8sgQpun
TzZrdy86k2uojdvieQoeKT0fbESUAmRmEHqbLaTDpKQGMEr1r3aUKkKxqZmIl7SMmtawLujE696m
OhSuk4dI4n2GUlMLipTClPoCHCasBcV8v/2t/Np+lxMEAvENQmu4zfj2RT0kIbAADikR7jIHFx3b
AdXciQSn3js85a3XMHdiXLFRE73EB5Rcj9uu1HBqgvaG5oHwuuXnJpDgIUUhN9g/MkBq8Yuyn3iK
eJgsWOrY4rujOt6hEXc2q21qD8/uoOSoBpkT5n2Va39LOs/a0LvqSoRo81RrxAftFiCUSXNCtTO3
+SRxrKSF3D8oWC+CoWUAH8iQcTV1HJeuRwNNTn9ANi3F3IFy2BPKpPcfe12wNg/2FVXcdS+F4v/3
2HqzT6x+ppYXgWpqoqXonTASKnLPGyYZJCACiqXIqUhdLtfwMDdkKpBw9PUYVEV8cG2KXUjtIdF7
vFN26KmQKvrzkNHl/BPYreev1RgBPA1wC8c3HhRrsVZTWQHjr+fX7Tq0igXmKA7+9TAY16MuTEu2
l61iPkpuE5WEY2Fz4YN7CtNV72x/F63fj3lGHmuBByvWpcOVDLD1/E1zCeiRy6vquawQTD0RbAVW
4BsyoF/AKp0H16Qa39wC6UH2f8PH5kJZeMhvK144JjLV5p2KpGmCC2/TVH1EZLZexZ9aWcXXpT0N
O3eeYdGokN+QVbM1GOrJoFIT67K/O8hyqTYcdH4j6uESlcTNHV4Hu61p+tfRu3byx+WAvA6waeeS
JeLep4WvGGv4FMPXiYyv8n/NsWouTfl8Rj4yM7Smn8v8HSweK3WZW4kJKcAI6FP+4U4oUASJmWWv
T2Rx5hgjsZuLmaUj2BZXCQA/qz2F/rSBL28XiYwfVYy55Vwqxdm8fLUeSBtFJK1bxpb6xYv4J78W
1N09PqhJvmNXpibBzmCVwPBrjhrHMIP2W9wv1rHttft+X6KHKg3xlI8AqjsIs2dSJCbpdniZlbMr
GpJGnEBdzJWXGmPcY2dRAeXfsiy71zhVcQAY2veeb2n8SwdwKxdhKYRsPTJ5uVP/ev3cUiAlF+sT
kuQJkYkNBzcXUR8+veImvWZB7rOfrQeQ2NeYgyBqCbj/ANUAXLEOv+kp8Bw1yKHCS1NSPWdDQhZu
EVATA8QYKaexzgrSn4tkce0B02QymK1QQhbkSbYDpE05x/i5M95xYWKz4hwIFHAlDxsqlboWD3A/
YQxffMf3f9v341WuHMY7lcaiytdZ9vNVAU5T42A7/XNRm/3jnsEHb+H326CNvhtfsc7tJFc+88gM
fcUKPdlPMEEVfJ2Kq94hUJCR1YcdrmfLwQ9AqYOWsLSjgqWo6Yis8GCl5++P570pgf3lWeAnnNRn
u0tN42X7SB86ip3dbOBbNBApFf8zHVFy7C1FtQnJ7zpiMj8//p6ucNHbu8Dr0CfmgnFqreuTnpfW
cQ5stvG69Ys4J4SH0UViaRA6iVSvdlX6REippXQ6NhgeT84zD5uPPjy9U/PfBWkvZSO5XewW0Z3A
tK/yJHstw+MnddWY0ajddGgRRAbNBIkUaUyhjLAzVZiFBJfrONIGVC/U4l2A/nF+xkWMxj14dHb8
iAIlxdQU8yM1Lxnr6J4F2tb+mE+FNXrh8I9PZvC5qAekZsPGpChJDOs0+3Rk8yB6s6fTbnOtxX5H
bilWlO2Fit4t3X+11uReGid/XIrZxcffLysaizjlmeBUofGiIN7o4GVZrrtFNXxbZocppCPu9nwZ
qxAmn0mMg9kAIvyIGnWaGks8FYYjhZmyUbQK6abmF6m/dGQFaEEAuARChrmUZVyU7gasKt4Zmp1y
hmXq7eLZYqujsvzNORsbPotTreYVRFWksihWoypmYDO7UNVh6mvHRHxZhvSTnhezODqE4xOLaAns
Se1tzs5JeQXpbgytki/1sRrcT3vZzneVtXJVpcGt6Eg4PTy4ns+H0ZfNrh2OAAK2LBcNUw2c+Mqu
XhKAz7SsE8ALBf+sKcx+EBfH+3aqhzNzDr3yGCBUE6IXnW+OQPtpT4ST+hKNyd3Whn0MilqrDmJh
B8Ai0isgqHYkw6DNBHhsKBDVw0DSDyU6p61XKi26+Df2r4DVVmv4VNuCYRDd4gWM/OuhQssUWWPS
LndBl1Sy1p4ApWVGMD+kIN1US/mlBGsiYYC/2sPoJQLVqkGNrdW77BBNmYNc70WZYynhaL/LSAUP
j0RFA30Q4+yCaRG+1LbX+1BcGLUzXODrTD9ffk7+PdnSHe54fyUPHCRP9Hz9O26eSgxr86sF6BDE
SI2jyGRzTCI0NSE8ElhXKrISlt0r4MoHVsNFN6VVMi+eeIHnxwp7jDtO1cZrHh9A3Y8Ut1X3SGBp
7QTF2kuc+dlYENDtdR+mbbOi3HJ6ax9AS0KdLyLRQx8I/7WlHgJgHQMOSRvbyeS1TzTOYTPEerwF
AEnzKfm6btRWKuXZsthAEzYjJ8JMRy/cYZ9X1QlQT6cxO3a6q9g2RpkFDS6BL+ssLgexZRYGV8gL
ruata6FWzOdA66HWLW7CQgDgMhu5GVHvIkWYh8BvqcBGh8iRtcgDHa9NXD0Wh1v6et4JOaXeqJZV
kQmwsPXCT/vqB/OyKcpzti1wFQ0J250mlrklGJPDfppXXw8hHT0wjc0EAye7EtnzYPPf/4q7pKpj
POrmgF/iE2XX1bea/RbNaQTTFlmIL045nqPeuMZiVNiYuJr8jwTm/lrslsO5bUTKSX54ZqO3RXpQ
StzqqNx9WMm/kXPaUWwvgwatuY5zh3+SF6rvbZPoNlOT9z1b3ZERMYki6MQMX2ONCR6jWy1EnO1w
x3/iJuqJQTY8ntMhnPIjrf9HYEUaUxha5S0eAxt9/Ed+JmlYs6iLitDqkV476IJUloCFQN2Mhl/d
2TL6BDSQD+OgKIogXXX1jS4JJFQ5Zz8Hwzyx4Siz358wKEW601SEmVvuHiTRYyI0L95kLEbefQm7
quQDhQAugGtHIw62F0k3GDdkK2mpwUhb5+kHrTjJ5PleLrjRYPPuVesedCoA5AWSeTkxRiGU13DX
qFq7mZzPil9nVflrJd/jZ+IlmmEfGwYtz6oDwnTz//P52VAqyLSSgGYQpdcKkRfpX17gjGWuS01d
ePl2obHLLYZIqEbO+HbLVnkUvFimpceOb0/32ISnPcOlDPiWMnJFfxi6mazNJ9Mb29gW4JDY/MNA
fmDx8SjJeV3iAUPqpQPL+LrP/7o49vLQN7mssezJWvbKR1109+E8h1/uikIqgbP3ZuY3s3iRQpzV
kLQ1CkBRRrBtX5RaUB+EnnEVLyWUrargTJcIXGxLtbJfBhH4uv3L4JkGCyhuIjCYuWLICk/7YyGQ
BKTn/wWIXWMvOVx6oI6Znj4a+qnS/Fwvp7QvRtoECliTTjIk1MdRze4i6y6yzpxKMr5cDdM8Tcdf
LPra4vziL4CvK/0iBo6kwlhepE2YqaOwz1ow6EzoV6C/0cFT+mwse/ytar261aK1Fi4zB2YzeWgo
jNpXP5HFfLCNUanOT5vyaHL9xIbot9KuES/alo3Lh6X+fllxd4cXxnCzuBdgTEsBZEZxjTKMvl+d
QRlRqZQtlZCR2JqWcmch9L2WkyWBhUGkuCvznHi8Y8XHKhVbr17R/V249VenIsiaPBBWCSfFZ0J3
6PVKH7s4aItbvS5tHMzQrjdTlL88Hcn9bXkY2u2a/nClXcuGTY2WTp7l79H53VKsSqbNr/LiNBRR
VU5SjVrHyJt7EHO9jVp3VaWaGRXI/OGiyvmUhIn+xngAyvvX06WdmEw2o1VfRkJsQzdV+somxbGd
/EasGh1WLmp5OOqJRikzH3CyxqkP8wNT3WdFtYtbApebqSdYQMkHBYlgqw8+b/4DPaJwvP5nC7hQ
lImkoSjsnhVyTfMeCfueA0sXgSrz1fq4OmZgs1h00t/R6r5F5Na8t5CPCjsTCqlxuTQ8tFVdTZb6
2MF0E6AtdhIeVtDy2KngT5F3ZQ3Zeg75bqLR+3A5ADm0G+F+JZSeEWuY7UuyMHk3gCmCnj7g/Nv3
HLUJlMx6qz7hURLBYq6iwQeqfNpWwpCTWES/FrR2sqKharyInLnoqDs4RWjKunNpeQxYVxV7YY9U
ZvFPI9cbV1FXfZHdLsjIO+IjXVNUrB+dR0O8MdVGHtaJKqigGBjaYhGRvrk154PcNXVEeq0z+D++
1LI+YJB2k69064CAXaNLA1AHZ9hQ+NAo+1Sg1QVWwxhrlBpf754ibGrAtCSvtJHt+8hK83HoZn0y
E3pBMuQTl40xrLvcc1nmPXpW65rgGSQ1HBbyzs9AIJ5mHVL7OrilClznuC3vEOST5lesBTWQ7wtE
S1DNmYBB/+gOY/J0moGQ60BmD0oIm5XJHEVRU1bQDNXvE9yydyWOC+C3NFizxdavdYbpvVPKC92h
yA/W27l7eaeDwYpEcSoALy7oIbrFdk1lz/kcpp4ISyt1RTwDUsD2oLtd9AjMcLtJw+pmiOhL/j66
x+j2KrhFEbdsUGBOhkcQ8/rWXGySmEn5tn+YspcnlhBQLLAkg9j86T89ijrJFdRVVHiZRiFkYUDK
iF88VQz7nD3W5XYeY2FpTJA2pu60+B4pYtSBlpIJrJLhULCqlOjJH6hJJUYVq15G3JD3mVDZRnEu
Wk9S+oghEiAx7K0RZc7SM/RRZemtjLwYjGTrDlOnQFEreFTnDjGSkDA1f1dKi73iKNut4u8s6pZy
b/xvIKHs4DsIPuNHU49p0q/Bz6r0qiX6eT/6fIkfFPJC/zM7uaubO79mRGEvh3XXyX2/dhbXm27r
UnvtGQgeYebIcxByLpUN5mnCz6030UGbmGR24LILt0VIOS6aAB9zxeMZm0SNKjqpaqQ6LP/0doe2
F79oh+hStbBDK3p2mpxnA/gKwDu/xbN8MCuNWB1W7hE5ENHmCVE3GQoOWhfONZfUQ+r+yqRaxzE6
/Pc14M2Y5hmyO7sKIMXOjyYb1uaQVFpqxE4I4Tn2LYsm79MbMSl0BJj3OzUax6obFeR0Vxz4jE36
yQiObyoJ5XQJz+VBd6C21hldAgoeyQo8VQAcznOUt3iBb/4YimlsF9dBTB6Ls6ETjhBtObAcVU1t
MA0ztT9P15cjfuhGhR2biFBrNiV+g1ZTJD5aCm4XEmdkPcsxHdiYkAY6S72BeQoxWhcuBCPkpDAX
KrSp4XSlTpD27zOm6IWfQZDdU07nqF+7b2+5LZZ7MkFqcsxCJ17TYbcuKrYmwLrc7xgJtun86Qat
fKieYnKEX4Yga38Me7lCqiLAWUY4IetYXvD8RizKoUZM3aOVZW7SQJFMepdJR3rufhqL3kb/zkAh
f+qEfsJCZ+JZ68C97nQeRYpmqLLUWOkVJEocRQYCtePr0S855WwwGmevVUSHNgFpi0SdFgBaZl89
B3teWcwfFexWjpbO6Vb2h7PIg8L2IDq26DKa+7n0Xcso655lj+CURUCPh/7NkfwlPl2HkCApPg+j
hgPnD41e4fXbfl9yBzX0Js1+OdH1HebNtsKwseHxVptehCOQVHI5pV/rSKS8Fm/8Cd4BBr9QEU5S
FVqgQVEPlNoh2LUQE461wk/dyR4YBNFDbLsm0ti7d0B7Qw3eDU/zQaW+wesNxMlLf0C6iPVqtGl7
VhKIuZNrcO/jL6FlgkNVRkp6aGCaa7JoLZVMBf+R40mjQ9YAo8tQL42HXwWeDVqSR8C5GSOav8jA
ytg6cuRnNx5O0oCU0IbYxiRvtZid1hLOkrZdyC3gbbcet2QLwKu/bAbuTxrC6LiXpfho2pu9Y/Ak
oLIule0wuUmUfoiCFaMA7xTFa18c+OB+pqC+EQ9xa9GnjdIBTuHVlz/pGKreN6uk5FCbLFCTZDry
zK/OaO9K7WF0XhU/21kCAy5sMGjlvH9Jx7ZOQuXsrUBvKg4RlVikccnThKstdBjwTETl0ZL9ozU+
xOwQ+cRS8+ZtpdMC4M+8eVWNx35ACtXvmu3RCYwsPKeE8p9kXE5+ddFL+P7u0ZikeORloy/sx1b8
b+C7Scf/HZRtM5kBBFDrYo8VoX0owqb0ODxpcSewlyIXXxhtzhVG5xlRY0/4+SQHuu1nW/YiCT3I
oZBo9/e4x0UnxHJnyRfx30Xkq/nHzDhDLFKBiNpnO0qfgled3fVL7XamPaXkb6J9WZe8t5nNHYgK
F9tlj7GbWJ4wBONZkSclio0hJUQNdJkbgwrRLAln1Mj9OkUE+VhpDxuAgJmA28XK7yYDtec7yZG8
ksf4x4L1PFvPgMtOMLePc4t/Yzp2ggXiQT58ZURI0wqFz6vjFwLbK6N6OBBro2Gx7+YlL/848Ano
TKQljFPMgZLuRhyEceddMqAq0Ddf1O8ee/rry6C98rK/9Onwx7Xt17OB65uPkPJfXPU9bKBxutAM
Ynp5xIOVLu4gnrQqGKnnu5pbAG1b7OQGNPsD2LK+Amrg9PclcwfVyV9uZ4s9xW2sZnizp7ItsU0q
ItVwEb8pxLpYCsPsOeV0MyuXQgP9EyqKSEPLhZ8NUVf6kLBgnDKykUIBuaYX5yPsDewbtxrwl3dY
G1EtGhqXxbbZ9e0NsZuXIIbMZu/N8nbCX6hX88OavM7SWbNr2hA3vordI9R3LV2ggcAf/9aR74Up
m3GWuewJPAw2WegwAJvxi06YvnTq6fGS93ngOEE6VZweF4R+Raj8zgMr2+TmnLgDhRtlPNnQ7ssM
KGMH6p2UAyRKcOpgXx+q26oCM0NZJJJrgoUSNiPaO5JaSIWNZrVuHEPH39tJeTuKcXzR6L0uoUi9
aQZJDr44ZaewJv8a1Wu8UhUA0ys4UBj952c64+s05OYXeSqfZSIadSmT5dRzEv5a6liEzdUY9BqE
WM6HmF7Gx0zd8XFdRoz0nuJeKoa1PmFBSNZL33QHTAdxv/7+qBTafDwyFWaPmrHB4uZBfIu+0YUW
Ab3jLvjasAEPME38AXc9wFT9oUtYHhi/+bap2JBxy0sv0G8fpzhzqJYC3gck/fjDmvizwoU8WBx8
N1fhEbl02MGXOf70UYTJPbIbFY5VO/SmqOgZGkekynCaVv2FiQyBqtJaQrvkImXg+8nJe/6JUFVQ
SmbtqBc/AmVYrApM4cKhkXK8xHspjMr4b1qOiz/Al4y/DglUqOFAuZwBdqnq9gS4gkajrwsA3oN6
ye5QLGV7dCkCrYRH/D36uWiuRN9cppSNaDx+gHhmAZgadThdwHLTfOsjglZ8KVwr9ER8Uv3wMk/o
rVkcToCU9x75qk/wplJxgAm0Z/u8U2Qo85quY5bHQIu4w4T51lgJpYYiYpOFqakpWFTYMwlR4Cab
dJ53aVwOT4jzwKSa5g21dl3PJWEp+pUturcVtGsXQADGau4ZhLjKUpTfcOKCH19LMA9thLY0GR7W
uelWU01ZjKPp1T6PnHpcryZLZsSEUxe7QFtuARQvokG7j3r9W9HBA7kNnGrEL6odostB6oHe+Ga7
+KfreFDc+sTgk2jMoU7LlCVsIL/G+bb5ow4xCkRrRdv/+Izrig9HiaP3Mht1vN8+KIN5MgEiFJ+7
P2x2WoNezwNDpgVBWinnjWOOO8jQpxF/BovOa9O5zuNgvdsbALsdgHShgKYjTnwQTCJ8iv6zQson
9P4abHy50UGWfXzzDsjyAknu+zbctdGF/oKq7u6h3m5tT5N6LZ2ep9jAVH0Vcrzlku9/N6LEit0P
vkuplKB9KvyN9cbY58rC0ni+VD7HYWD/0QTlkir2MBWi9tEC9M1JY77xNrH53DLWRg9HPjNoHI6F
IVDaMhKZS8o7830sazgYv+89wJQNzlnaxKafi8kao67g7EOBy4aSBhBBOmYFZEiIBq2w+EpK9sRV
HIlD5HxXQeFbUtxdf9fWktN6+NV5eDMjsJZo9O+9MeX99luFKe4rGDb0uxf03ThdWM+pVv12SNDD
XPlTPv3aVhfg7uLJPuG6ieXPuObtjwENSxf+oeOXK25vMD0naZxdgtHXF5uBlyNaMohQ0tR7kt6f
lltcWP83tzco6NT3MR5gV25LpcJXrKViOMyzhp7lhIUwjRn398elCp3KJguQps+BbtvylANCklEx
82tq1If+4yDsPAgUCRe73M13Kvm12AGPslOL09+IImc0u+m3VUzV1epdBdtKEe9EfvSazCuTiLij
XIkNWRxOofL83Q/6vQAxjYxqydpdvouS40G2Ac5OHo618hO1r5GrYs56ePA6EGkX8BMLOrdAQvmK
oH5N6/MjA3ImFVAVLUKilY+aEjHXVzHcxTcmGcjebOJBmus+nsvdWYADoQEyURHXW7hXYNvvthiA
elFDid2a68aGEjdJjh2oHQ0AtlEg+wkyLHNPCa7/oEbltxfu0yYtsxXtunhBuqg1/sMN5tny/a3g
oLdkLTptsl6yFbRoC8p+ZAbQrQ+iQnwb43hDhKIs7kWVouAE9ptNLxPTGBFcTXbR5pdF1E6o+oKs
1HaqmTjCeUfpEJoKEYhLW99DW4YVxTa9e8cBjrsMtDCrgwNTs7XYAMK5zU4yBGKDMvbVyTE0WXuw
aIMPnySDgGk/s0jqrtPHgLIigHEPJTAeY7je5sWpYe9xFvgGrqHewkRa+6P1s70vbK5YazTne/nD
7FKJwKyKpbjdO3Gy83D9VHPGDM1b+KfhXFbzPGiI/+as1HEIoAHGL0O2ByH8HGNpoK5oJ68IZx99
ODVAvsyYAp4CUoPrEZVwEsVoxjUHz703dViolMG7J3gkjYlT4IMUk9/aPxdSa+2I49TAc5bkK7Af
Nj9+cn6/fGi2T42cnvzugfWKWQtnFnnyuvVE6/yP7rxp1CzK1Ukc3BAAjo9VouJwTY+e/wGTihxO
tVPQ4PgQ8E0TWPuhXu04hHZ3IYuX4Yi4q0XwKvJTSF4PXbaPaqy0bzuG6K8YVc3ZYyuofNRPVc1T
paTzAOf6J2mcYm2JqZijXZFkiJyo5VUYCsORnkT6ru1/P/TzJCkmH+U5gRe049f6OQ2f/rWZk4dr
s5zKpez+Lj81GAh6qFNK973UA/M2nQHIbyrVz7zIifRZTsXv7WNb6QB9lJz84ld5/DU5E4bTQ2WA
0V5i7I0QsNqjoBW71IMjB9xO2K+8u7ecgNCWj1eJ2c5UC52UwpwuxxZE5QK/N844OpZ87P/88GC6
JDTxV+pRenXxwgfneD6opbnFUqm/X4iMc3OGGwztHE6ISdsPn1lCyrP8v4/GS4pkjkLqNI4ns+qg
4LwyptD86c1noB1a7/QVj3ApkFeEKV0PUN+opunA/wLmYUfCpnNilP3FswKEPZwYju3PadLuboPW
Dc5mJgf89YSTaIcbXNHiok0gv/Q/jtHoR9pcktyQDStIw6Dcmfy05KPexOhKOIuTHNHofDSaB0A8
dLxHjZgjBL4rly5g4PBvJ2++dINne6GgHGdZmrXc0dIHEpssdXWZ/xsR7qBeovCAb99YHq5Zynwl
qPvFyBOFmSEUNCt0CzHrWQAimHeM3amRU4EDiuzZC9kI45ocUAd9/Qe6fVLTBZIg0tx3Xfu/PZDL
9/BOTggCGhJeOxtEchNyCvapywNxeG4ASQ9CUL+HuqmGjUeFqt5elIJJBHPhwJ+TjTEB3qhzrt8A
HpjUU8Ev9PuVyTJa/Wpq+tvMLr85E00cHMGbizLPLwf473KndwvE1vOC532754RkyWf6alHFnG2l
bUOIV4ga+kVAi90UYiaDuIZjHICpW/H0cX+5lPQ/0FIusVJwT9IzNJXKBzt1K2BdtfHzWdE0piiO
8wacTSUFdPyxv3p6gFbMbRXXuEntlUB9On7HqrsrCzx1Hfo+C/c1TF4ACzyv0lxVEU3g+LHv4y7J
NcTdSkL5NJ2v0nma2blUODBrjzFXbTLix57Ovk9CRqYKUu5PanbNznfsJycH1B6C2ENfj6XeyzqF
KcRSryKUrwut8ukjOMeXZsRJpsdT3zlcuWCYOsHmHnDKEjkKk/UmaPam5CSpbgIl8j+GExwSnlZK
tEw9yqt/j9yhD8VRgtjnV2o+7EkemUrbehvTNnn8AxSNsUbAnb5g5/3x5su/DkMFrdUR10qpe4Ep
b9kyrQTdNLXSGRQzIWDy023GbCEOEkwJ65bqgot7ZwQgzZvLL3+8e4ZBtZUcpVKNN7DLsI18PCDS
ul1dchJe9bep6DglZ1tgOnDH8DwjtBpOzEtQvtnML08+LRWRMARrtWDKpiFWzBwU5S9DIFlJx/WC
lW479ZCEnMcLArrVvl9HE6ZqpWV6QebxmaE4A78vJd1nH6UCQ6m4borvzehECah2VSUbuRdqMY/g
J1wmPXUC5SOLlLZnnXzVpjzfbN+AC7qN3iQw/gWGGtA5KTiSvnaHKDQLYsFmMq/1hCpgjmKhmQMx
hT33qFvS9mbWwkB2H22yjXKKUFtiPQO8go2Ec3X1s73pb0FYP7yi7EfxQmm4ikNB7aOu8pPgfPPQ
niP8HzabeK3ZU5/kOSQxYHQenQWjbz5iWME4U5NUUxxmjNDYXek6LMXn22F41b3STOaUphoPOXjA
5Wl288iDWMFh0Yn3tiKtDu9rB+oIkqhUPOEAYgf5Ut4ghsaZvIAFjeC/UueovZ4wtaUY+w7+joti
rp4paFPR87mRAD+tkDK0KYCu4IsmI945XovJkxLBko1lk2vEeBCuyL5zcQQEiQEj1f3As2waiAtk
CCLUcy9hmfwLfDURiU9jKm4JXqIIK/3CptDS32tjClvsBt9k//3coOJGWAJKmFgMYgxIgtYTUmtV
eytShAamr+y4N40dYFgYlYBI+ZoOxK2PqStrWwvOID9s4pruBB+Fa40OKe4aaAH6NWE8kDKve9wT
RvgbhizQ41qeQB0WXd2sWgI6HC+3rh63luYTOqNupo4w9HJUoqZ3VGXRNHLRaRi8/otn5qqtyTZF
Kkm9Gpek3Jo8gzLXwiicfTLYjFu8UfIHKCrCR080TngMXZx5qPfN+jJs66hTpG6RyIVnnx8uqf20
Tq7CtWR1eBBTMqH2TlO4HR9fqwgYEkghy3upX+/AyV8/I4E9OxZiUThy1kc0ncx4MgHyiN+Vbstj
AE86aJ/DzIy1JVPIUkvI3MxO+u0qDUwLKe6U21bnzJz6jJQ56hsWWFN7zzlsHUdji4AQmXOhAwHv
oSqpDs517YOjbTaDs7e4TsQ1k5pDikCXrDf6DoQ5k6fdRg+jd3f1jLCjYxPFi2vVG9AQiq+523r+
Wc8O6xdIvH6zv7l6xQW+ogj8jibplQPleCrvBZjGR+vE6YxIuI4oOs9/5v8uOouJk/me5GJnlM3+
DiRLMxFa8aZMXnOrMB0z6fi2GFERY0oXKIW3WvKSnRCisUFKpABbQu9pRDjqgQbH2mHEKSY5uK+Q
56ATe9r4zJ+xdE5PJA+68DtjvNXs1d6LDf799C7JdN2b5s44SoS070FbLNuVkm8EG45LyDBiYAVs
UngxTmGxtC0RYZB0/Fm+qb2HUW5GMGbWIdqQYxqZhCOVy1NvVCrYI9uexl0ZyAYgoFcub/gGsH/G
XkyWJN95ECdqfBBvsu+mn1b8+epabVss1wj3QzSEkeYoq5XA0DmFLqqvFNYXtkWK/dStzBcrRucn
2nulfLHQS4FezViuHx7tPVwBCzNLqY8FRFIsJoOWuU+xFfIw4xATu1Ic4RBldtdrrAo5Oj75Q9WV
BkyworWZrXxtYkYNm9xRnHyVS567vg9r4NgiRGf/gQ5QOF4jKERvTdMQw8cEbjTSe5BV0oMfrJEo
IgDO0A4CG6wiBG/TpL494e/myh9byHxqjuLmSqua9G+CxRAL5Rb8+tQBc5+IgXRsD8of+pNxjaMy
a4K1GMpTY7kLYK1j98Y79dN/2VMZT9pINEU38Q+uoDMBzJsDHj3AR+elwB88oGUa2SELEY+Rcq8/
fctaEuq3lnc/xPLCM0RIGaW3kN+9XV4tqU2p0AwnfP7m6yjSIkI7aFaAYruqAX9TLhfyef9nAK4d
0pfIXXR0Y1CId5X57wE4uHQ14DoL5n36rOTPNQwHrHn8ji4UXHdzw8WLYOuRR8ZlxIhhU/52gnDX
WNcax1WlkisSjVTeMJjOwa3iTwIEv564hxw0nnALLdJ613Y61uqGma7twGKdFOsoq4jLR/PciAtu
GeJk+Q9ve5tujuqRX3kIdgWB4LzBo1D2zk3WCFTv9jDFqGEAmixJYXmy0SA5N5BzVKT6/j1jIIUD
k1TuJgAqaDe1hyRz9De11oEeTdIPmikEUZQMgLUBPD6F9Urt8tBErD1kNxGEUnbtrrA81/62Wn8Q
xdDhF1SLaKDuTkwXeGxJptL0v4yZdK/Z4cEl+dIT9mlW5/N5j5rOkmijoP8fnEsMe7dkPyCnPz66
1q8rAuaCtPuMlG+RvqqiGH9GgJXQEIoillwxvls1yPDemubX/Vl90Gki/3ksJBuJzWn7rPjBqAFK
2jXgzzJyKQrf65q+8FoEUnwWiSovthR0nQgObHqLSdNtpB8LdlXXTcZmxkn/j4CMz7Ru938YJnrA
t+9XXY0Aeq7VZan1vVM29JyxB0K/ixQ9lXQpG5ts80JQrpfjfjh26Ra7ahiA/ha53ZC1z02KXuiv
mMpyApZg6uRZp9iSCL2CTmGLAFFS5/bivuX4Gr/cPiWHuzAx5cMN+i2qasG+YVdnb7YhbRVSVyKo
4Ysib8arBlOmd9jdMEEn0thfX61H5kNIW7ld6dskwAg46U8DYdDFeV4lJnyIYlIPrx3CYxpyIWO1
CQxTFAenMZaWDjxPN4C4y0AtiC3SkK+os3bD8x0DUEUcfGsn81ou5xZ9/QxbE8JmYWK4R4/DyGYt
RArxj7zOEwMtWzaXWoioTCNqVwyVpQ8bRh3PslCnUKhyT1Rh/j6/VaG+fO7JfeFaI27SxLdFgRUk
eNbTfLlI2Fx5OM6u0LTWa12AyV6vDVDoVDygg4Cmqkl+P//W6DTMlXwdbRY6l//UGMvs6x+SCjx2
MgLzQyZRnvYs1t/aWLPEfSf0wmtp6tRgW5vhaTKVxn6NmHTHfe+NQkDkUlbX6EA0GpT4Df1STHNa
zSwNPAKj2L2lbue2d1QRXxvRsiLUL1WG7x0JDTlYUxtT2sFb3yS6WQObXZq13zygZQvK1F8EJF8C
kf/Mr9toZ/61bJVulHEzdElJnyVSwBAo2X8guyU6qszS7WI+oD0IOIfzC3disg+qS8QMezA8/2LG
Xofa6KeNW/aacR8eGXkPAWad5V31ZO2ay+eH9Uaqo3YSYqfZ+F14ZHp/MQwOcZGhQuZHEcI4UI83
5BONfwHLGl6plUrItNSUJwpsvpoSVACrzRFQq/ffI7qan3Ur8PycfH3Ya0sSURlZbPmHfIwnsu/3
fzmCdnwrhj+9XdzH3RRlgAJSWuM84uSO7u/7Bp3cBgGZH6fbFYlIFVBT0N7I1AbMJCnudjl+Jgv+
Mr8g1ZlARaszdkZ11llqMUWYdyYYbqIAGry6b9ljytP2Wtv9G5Z8o2vhxjn/m2jTKYc4e9QYKnad
E3+us9UBckE4BpRA6dBU0/ALyOWyXSC4lhMOkxAK61JrlfVnHEb+i2XCVELBGClfgsYehFsDgoVK
nJ4Cefvwgpg6zYItkEPvmfNmlmxyiS5s8cEQY6QrUzCOO3/1GRW1lZmR3L0nCumvCxoRK/ywwQvi
ag0zqUbLg6SQXtpHRLRplJbFGfmFZBRlP3KjBE7dpn5W8xJm+TZ0nbvr/Cqel10gAUVBurvYbcR/
KKP+sPA5QMJqvP9eEPIxQdkrXQvkwjFg1L/agWxGfkgiCZCWjmVRNTAsHeqLn1ltNfGTQK7paqKh
FLMD0s6S3L3wRxSQoyeAykJzUSybXXSs9XZmdSqI+NMpANpPO2AGv2cUSTpPTnoUi5G70/6VnxPs
iWYF9IvaoEYOHFibxemV+BJBrAvVeytRwcYgkTRp7citDFIi38vFTlKLFo1zTnaJd6XyzBedTNao
tHXBU9d4BATE6JDwVQQI9VbWZelLL98wUhePnaE8xTSNGpkJ/VYFVRrIrMz0IBCtFDerQ+mS9o9D
TkjOJefZbZiqfUdmJ3Vas0gMh05Yy9TjuiHQHWNguMh0FsAI4rjB+NdBUmQNAvyVE1SD671p2fyh
PL/aSzliTwepUX3revdKZaXjSrHx7bqzNReq+IFPyG6c1oQpGlyaNHpC1FgFEAjdW4bzR4ixJVai
fzbQXAeWYJiuJb8/GLUUR1b2zFVu0XezDB/BIuJIL+RgtvHHde+WC2TxHR6WBrF2MBnyGoatHADQ
r1QwbL82SWRBosqiawTgS8LCucGfdrwR0uh2wE+Q1VFt4BhKwrQhdj33VhdkPxxfY5JBvcO7Knt3
h4ms9AUF7LQPkMBm1VvheREVAvts3JgmbeZhAc4H1WUPDU6J/U5XYyf72NgmDZytZRqDiVvfUFwC
xN+5xo11e+UYGHjxkCf/qkahX+LC5NTnIOui9IZKw8Ozd32pChpizQqsF1Ys9GYx7+JnXghKz4w3
GczyV7LRcukxp6/I2bIyVrPFz4XTCiUyc2Lr24eeCjvikVAQRSdVyNFQ+4SVMG40QDNeabNQeai6
lxQChkGRIDIqEl4oEg00cFtAE5EAbhcghHR4MucVSlz7YIXvZUzluiSJbRAQe3xN3fg5d0aLfMqZ
Zz09Yuz/pCeqyF4ABjFjUSSMk1q5b0Pv/jDh3gr03RMqcoNoguF41XrPYUIUDXz0wpQnJcM3nuJd
6FR2uQ3YzTeG6gwyzA2mHpQ3U+wfH8QlHOhST2o/q7tIUd2FZze+s040ytkiaAwcRwIVcybrp0QS
aQl9Y2/iPSOnSYqU1UZ5rZRMnuVTVIZqyqytxurzO3Qe6Nu/a51mRxhKthz8WIBKtQAuTJ8aMJjq
Wh3Cm7c/sb4N/6l3Wu2yW0KTHQB8yHSfomED65UR0gbaeQTNkZZkykLPjB77tEPtOBXS/fCJE2R4
CkOFyQ7QA24UdgOlqilouRAkCZgAQMxUpGSVjo2gi4F1kyzzeb4vjeJN/x+wE4zQHm85VoxJNZiv
nK+1r9wNs+8Q9TKmGx3Y7j11fR+rLa7K/MDHMpEMYxszcc6JuTLOTaz/bRBZxdSx4JnpWWJhvb0x
xsTywSO6hv84ashQzN+fUzpXu8ckAU8Wbgml4GjzcuIW2mW5YO7rtrf3SvZrNhSfbhBmrf+UejLh
KRXJ85nR1D4SldHNNTXnHm4NtVgJWoS8JFS8C1P5bkbYZAAcx/u/YtFKICqZGTR4GQp6nkPfzu8a
ywtRokcTLBqdhL3mj6Xk/9FhMCZoZ7wrKq6qEXrXQtoG3pszk1X4H9bn59nnhav+C4x+IXHyOf8e
8tKXb55a03+r10BPjysEfTTVkw3GCUDU2avNWH0ST2/MIerYB92nJ3CpIifSAJ/nem2ivvox5HJM
glTxglBZ79jWsHjbiA3JPRbiMXBLd1Y/acUE0aurMIeCygZQY4QK/ONufImntQcLjOjfZSjW9qgI
VZx7t2wiGl7Bry2uscncpQGj39PH8l0ke8UB1jGh9eh1exmBR8yKDutz++aPk5cpz7aWdw/20QPa
oQvirBk0renAO4AwZ2Mo8aVQhcoqkBFm0W4GT2uUbkbQTmexzb4P1CpShapYPzkGNyWDeVPbGjGb
O9YXnfs8p2m7g88M4F0bDqNm1T78ep+GmF3uLRrVsOoG6x1fw2jriPEERstW/wbQePtaCLPa5dS+
2M34JvqUtbcKrHaj2H2KyUh+YFYOP3dANCjVSgDBCVltX+6DY+QG0+Ymf/RKpPCmqOKE6FR4GAhS
ssx4ex5QwkIm2b7QQ9IIMIxVAZykwOcDZY9LHM6ASIz6LdOJgeCcU+K2eu4f/qYr13F9kj7Mvt0W
VfG+rzwSNJ5rZdmtWg4YxRWf13Dwz5tX/LjG+WUpCz3YMXNVm4ekyVXG3N3zGEOZpq3HuuXJW+xp
Y8udn9A4PVClttHY/jIvNi6yPTK1o3jaJNfauQl9q/3mme3zN36AW2XVXRTC2Y4ppYKtfP9UlLAQ
FwweDVzvpQOJgDk/1aLu4N6jB8biLOMY0eV8L2VH3+Ef33X/0FPbZqclJMB8QtM2N430bkh/Fsnz
6BxvDj2N3ASeVSwRjUxtCmeehQFjykkP5wsH18mXGNC+a0RO7p2N/FYQH7cTkDM4R0Ywwkz0ZJ9l
qZRNjZ7mt8pq8di3sDkW2xuzq5uZ60CBznqvi9lG7pNztQujJtRaEmKEbJI9SKblWGJDW2EgBpEW
ZgglzWzovv9I/1iWVweEtF7xjD5Jy+R2i5lE2McQjU1DCFgKvBuYaILIaiHvRRbCq89KaQaWn5gn
sUfLjGuYCNe24PqEWlB8ZTbpCplvTsYeNnFNv5GGw538Jclm0q6qOh8mJRO8TeL3Fyy76OTiamwr
34YkumfSx9IpxsCdcz8PpKNvWqfFL9aNW/y8kYwPUenGKwGmFq+emhkDAQA5zz6ofoToTmmWrdfy
OR9lqXU2YsYJFPpI1noeaj/z0xg1n+IkJ/zb1O+vemBnCoGMAn3wNds7V8lHjAv42lFWTJeSvteO
1d2FFvnLMgo/o9aCj1VyvD9BT24loxsxqaQ+DKFah9mNfIiSPan8vnoIqp8QPwg/LbBseyTnJAmb
ujZm5ZFuebnC15WlxAyOCDgozk3UICziCfuv3E7X1okSLQGhek7+hi1W8EngXD/cip8QbS//RMJL
NbWspHFt4V5wvFSLkwSilsuN38MZClad5g5gIRslCHBuH70fv2jiRbIW48u43JolCMgGAyRCScIY
+HT2ulBzLImTVddt8cuyA+GM+2xsrfdXiKNSwZQyyuZ3+1eji4FR9pIpLgwH4vUl0G44SRUfT50d
s3voEBVmr0wPmqPhiBG5e1Wwio+NHlMJWEL+SZTcSohM2L9bTEz0mjRZtI8cFz668Mero0I5hp1x
/a++21xf8Hed+5NubBFs+eM3pzWyS7WYjQ5b5CVWDEIrwjr/X1+t++PXMVQKL7wvg7jnCV9oDLM7
WsHU9u9d6poSGTRJZV/d9u2eKDpuiaVsrY6yHN/AXq4F6mpT1eDmo/fvyzFcuiVevTFIuaeqqiFz
IHhtqqMqIMMnFB4/EkcDMJYxqhLo/lPbP/PnX1767nCDBfliDX2xFsDQWF3cthTYnTASqdJkN3CZ
lwRNLfwA0MiMYTWeIsppLcj0Jkeg3tTZRIOj8Q1gyP1ewq7+N+QDqCgJWU1/Xo4ZqvI3irNiay87
QXa6L+Lb88KecmM/0iftLECIyKLVoqmv7ZqtFYXzt7Ejez1wjwZP7sYdWCuCtrHaNvHOb+aw6CV5
8eLpGlOkbmHmCu6W4P0noQJmzGdlQv5fiFBnaSx/B9OvjhsviotYobe7T59Z8MAIaEGIEfPLFaHR
vrPiwP05N+yglT7Vny7vV/8nk7zTNToUZvirhDlfK4jnKiGK3C9Z+sieFTifEn7GpoPWKcetaCSU
rqhED+4ShDwZFxN6oCzhcn8IGlS94eKHl+XJTE4hDJ/FzGh5FzVOjlt+iTx+ZJQWFth7HZ9bIuAX
Di821c8ef4rkBxFzIOW6elE0qM0wD8CI7cFpjRe2/M8T1/hwkcr88/+O/aAffXgjK4xre8Mw3W5k
KPS+IiTQS+mSRFl3vt/CSjnt2xAk/a5xBQxrr5wpbIRMaIC9KyWT/xCYWoWQyPNCymNXJ+1j4v/4
dLe/ZayurUDZZfshQDxIt2M4cJCaZO4FjSFFY916oyG/PDMQufuBwCJ8p27Z30vc5asS2iy5I1mQ
VvwQUTrZA3lwYvFOY9voRsEpLFol67AR3WH07Z8CBKXGmREAzp85qF257r6SvNwvZEkjeVrkzYo+
xGODIrYvHofn6dy4Qqd3q+ogX14boIbogWb0KG+v1U0cKGNnd7HRZzlUKnt7S7VbhFiYJXaTXYcu
JjIcDYz/Wl5bkPSFU/xTw4V+RTkBXv0sE/rvlHoJMiSOPRv+bmfyRjSHoCNdyUUDgSxisHIn6ZYm
nA7eUQck+TfrO6ku1BixcolrQob/bSHlasiR00WUti59Dr17V7cgiO6320QOsdAJpqq19NyCMqnR
4rA6PfolGl9yQiluAYE3+5pNs2AhOdtbQi8GW6NI/QVoRyAN9PyEZxxiklVZKrmVBjQvZ5HH8yA3
6AGN0m8vpaL8DiKYWCqTqufee62kTxHVMipn6zENVLa+2rgYogJb6RZlPyFf9k3VjAFIY6Z2ZYLW
r2MJ07O8RRk4SE/3oM3d+ajCV8PNaFRqUp6tET2xFK5X2x4HQnJQ01HcdZruP9b9U8QwZeG6ecaL
PEopybvJSFP/E5LjgpgtlfaC6FzJ/nRWGV5dEbhvHjRplYmQevhlwGvlLj1qc8WFxJ1ZWtepVfsq
y+/MiFIuXP8bf9x3s6/LkbBRoWIhxjb41UVmUQS8YBQtPaDLqqzDMATn2vVStWK+AGJaF+h5KLpA
AsLat8cJFCWOKOMhNq0YOFTVUshBzHOg9gQ0aY7LHOGxtZ9UMncFuYqNwzzwIPeTFHA/XHowi+2+
jX18+orUOAsBJCkAEZ694ca2ojWvWGreOrpNUks7M5kAForQDjWRSLummmffMt1x+y9VloTcts7D
K0CaqCvMSTn8XkiI1P49NyBJXdCmMEn0VFYSgFwQsb4NZaWWXGP7b/ILp5BoB5hKd4IxFBl5I0OZ
rTQTaltqMvgtqTzaX7y4iPgWL4Z8xT2WYPg4oEoqLrTOnCOTQpqxJF6QGkH1rZ+yjDuXkFd+R7+U
/TJNO3OZKA8+04RB15hWhz6ZYCnx7rxx3yfki7RW7ESJVX3IOO4fSzAgiUgbYas/4S2s+IW0vhjR
LcGkNBDujI4O3DfaiJLERBoHWHHGbXg1iMBs8yWWC9iPkx9KBPi4dzVkny5fpL8gf+YV9Oo6Uxu4
bXZFdpWt2SHE4iycOMD2Zyt0nFXckTbEViqcZiEWVUdAPOYjIQrXpH5Gj3rL2LkhsHg14p9+2xUB
1TpAyvMDzH0hV7FI0+AtTn/AFogJ4UXjN1Wlib9B95Q3zOJdVpVAn3PVrnR672BTrN4A2mySknVR
77l6RBEqWd3DJm7I+qG/VIE99uFtHphsL0T2VDUgouCYBctKEBLEEiechtyEgC3hEV5jw1TzD/Ey
5tCPk0Ok54VDWFy+W6qkSCiL5DaViCs2e4baSxPZJOoT6tIYckobxeyOrr8O5zyfahd7r830blxB
nn4HTrdSi1Lt1c99azp8dJHuVDzaCn0Q5I7bBIE/JIdcU5Q8VjCp7R8pLyMWgI57WumIx/+16tCs
p6GkRvLj8cAbN16Qj/iMxhFK8PQcBuk4LP5mhAKiwG4mK3zARLoNIoA3ALsvvaL8mj588nFlKswP
PoupD88mJjEPacGvMyF5dxAXyUXwEypLkcxTiuO+ec6DfPWwlQeMbf/9f1bNZzHQCOaSiQN4TiyT
l5MmxNshI/uKiTxieR5/PwAS3x9vtNYQmcn7aOzB3wekQTXhBkbOLLRNE+2pDpNy2U5cgscsXTha
XLukoM1PFFxd7m4JPUVtGaAg8ozDB+3VQVYopKVc/k2uukPaTtt+r+P5ZBRxnGjLdlC43eWM3m6f
dyujzCcqXc5++NT3hIQazBu+QvonSdw3zJVp0QdIvxpE+j/0/XIDDTe1MooYRXlGYAr9chGrVP4l
7tzUlGLBtpBG62LU8qEMoXXpA2omCpaRxuLjRGPDaXY7PsFUdXk1dlf3vRiANyv8ziZbYHFYadlm
NXyTlbaLl1N5If7U9GDy3+Ds5ivnX6sw2eb+gNlD/GrKnc72uc0OfZaGJGg+h1OkYA1iAmLRYzC7
gU+9FuWYVS85CmLtzKXpJ1MeH3T//PNrUBwDHWUX8UVZ9D8HoEB1Qbi5AntYUX9RQZODQzKi3vXH
w4fBQu1ISUsdSQu5r2V0lmnKdQxv/nnlzHKiuFxB7A7jbzCjIS+jsU9d1boX6KwDCOjAzK7u0zD6
WyMmidYpYxOO/0xKLe5s2Q1VA8bDOQFWVP5tykTxBlU6b9DAsmO9TnAKWElzmsmIQzVsIVUnO6Qd
+8k1I6vdIHSm6Jll2Ec0DDpHIxflTXGTf5NWikiPGb9OQ8N5FrxO2eZO2FFDNMy9pwhcOGCBGA1u
Vw1Wc0DmBJLaW/P3okT5gO2hCCCnR5eElpwmumRFvMXmLIAck6XehbKTPl9yTCnjoxYwJCSMrFH2
GY2dXESCLbxhQAOUzpqf++uD/gXqkg92AimCkFAvDtQI+HquLa5Jz8DMkA5oIi6Ee069MZJ7EoRc
ZKl0Lz3dYtthOHqHr6W8H1KOCA8vZq3hPrJn+vZ+mFGWQL2VwgMg1wK5K5lapIdap4kVpLGLBBNC
kF5HS4iXR1CZCigxBFcOCOqJK0NNPtLxii9WeubnLpnEnCK87Dxi4Kv4L5babzDEpUYWAWjAWZbI
mmW89HfMjvgX8OXgGcjc5fStSkS5RdqdiFzUItAo/utGZvMcQlgMRVFHTl6DDBOpqkEeAZvkiDIU
sLCabxHEnwTBkNU1iLrycJYHDPzkiIyrwQI3dpCJqMln0LExQaqWm1qCgtvsYO7aw+pxntmyeEOE
nHyfcGsrqRvEZez2q+pZIrIG0/ui9pl7SJ6d0XEftnIYKeuSB0F0nX9jJtNljq8RQc15gaMchYzW
B80NcccmoLVc3ui9jBWKxNReNhAKh9LGKAiYe4IdaNCkT39U32dtGRDcZk6X8c3PyvDD6zt16mC1
dQyfYeSWibwTrhLGZFX1t8VBSKQR/iSqfxN62oUp4YtGTMNP1UvyMkEqiuExJ/W/x95i8GbRh2JT
jKRHTWPw49UGzTk+Uj5WzmKdGlXzbYZdZbz96C7MGjxrQK1yw2r8nVzlLylugqFPd1jVbyhAs2E0
VjjULS1g74LGzPWVkAXok7N3vsQs9gVtZYPyZnIMP9pftcoFE13D7pBvYi9OHUcmwMvA9HKtinto
CE/QvJEnRRwVLyOHHD3QiuIe+j7oLPQ/TkREWj/JOauo/1UfwZNkc8G/57Fi118pt/dIvjh4e9Ud
Az5b/EG9BvwwEGDUgDvW88XcLETEFOcE6mjpylKNJoYF0GVR1aqs7U/HbQjWpTWiqb8v8qiAgf4T
7/L3GHOd9XLADfk13RfXkVxty1LfnkB70vxYQZssfXM75MHBzuodO78lxQjDqT7AE0gjVa5y2+xu
CX2jpkVX96hH7Y78f0Hx2hCcXqSUB+cTQmRzQ0groMT5QZXef9zGFwIfFYVITVJk39EVpcFxcsSy
rTRdXY5y36Wm6TalOe6uGmEcioLKsCsgTSM+bCjn+eKqjQnWKSGqvj8GcHjO/cLkba2P/alWCPh+
BvPyJFKt69N1OWbrH3CGYgytdHPJW/Iby132ufbMzPkfR4zYu9MfmMQTOx9Vj+j8iMs+F3C3I6Og
qeNFqKoEAX2aUflptRMnKQ7EXWk6vUYIzffCh8pO8FS/wV3Go+6l3UCUApXyAsuq2jXz+aWAqM+C
jSec+QndYtMWwNBRHB+ZPodSHQh6/i2RxbfdwKhP/CrIgitd3lcpaTu4WUWYHl90j6EPabuyEsP/
ZMWkVWsurHkv3/L9eo/vt3PTv+RMNySt6RwzGPzGp+4VXzLgHPB+/gu+DCEC5Q+u26syi3lYja4y
uApdHRJdlVZZcxV9nWLNbNHUkKLlEt/g1ZTuDDT+3GwpLeXH2GUt4l3s1nSvaPToYb+r7cdpfbhw
fzksstpfmBQ3a3doIGKOilxu0JjLjYtL4wfd7QIyVvyERk/vnUN8Als/alqBWqbe/xA3/DWWztfZ
UfRFV5a+LNXqXqp7UyKDBpUwOdc3nGSzH8/ZQ/FtXfFtWAve4SQjyDT4H7RVC2+SoOJq+9fQ75zC
5q+VxKPxToDUtu1pTHOiH3rXt4ArkUlKJ6mqkw09gcsFo24yiL8T1HX0biMncPrvcplGUS6Npbf/
cJmE4QJhpIANVlgm7coClnS3ipP9SrGOdmrJZgImk+PTAVTn1mjpvd50veKISw/aU6FbT0ECHbk9
zqHSK8G/ZgUlD/zSHvKAgEfjkDawcNpcnHoZmu+NrOyYf467zB3JNn7TyqhgQZA3OEHWFZLQY6eS
EMIluVMQ1WivxxZVGQPjNcKJgFFN6XkJkcCnTu3pJmwSLc4qa8voh/Uki6QtyXy6DBJlSv8OA1YS
QX3oHacW0JXRD1CPrc8qOMo4yPfYx6ISdSD8evWkmmRCqeLoukaDoWfFx8i2FEgyHwzlQ3kL99BA
mC+ETwUlDC6X6A+itqY4zL3HqGPx7DjE+PrJK7RrP5jkURPzaMOj/l59ne4d00CNbHnfkQEhtwUc
fsur4yRKFvG67MFhykMvkgq3Xx0eVKmoaeNzV78CiWvzoKt19cwRJdUAGwO2skrSTgBVf5xZhynW
lnw47hqLqaUnHNbt4GOwyVxGKBa+NOua7+XJu2RPYOA5fbfvvFBv1PTEWuQmu/Es+9weBoHb/PbM
DU2dupCoB9kEM2SUrOvvM8FltavlIA0LBeMIwOSaEtgFSvFycF3cbq1TE/57sGDRxPCR3PHhh/7A
oOhR/CVzyOLSQZlOD9n20wzvrOxly53XEhNvmpLRcw4qXEAb687hNI9ukwJsB2o4r2NREW3A3x2j
FQwntEi+GCSlD6BLl8JX8QZiKg8e3snsl8XgrUw+r0mT3ALYYR3vdlNMX+kPaR8eLbY/T48br4Jz
p6zDRYLDDhH2tI2Juffzy9sVjYKxzlcfygVCM1n0cvYDljFLgX6MjjhN97FYc5C0R8WmrF3Q8pE8
OSpo1cOXH6JaKK0aiPdDagMRkp1tZVYHrzrN89YjcMZzAPHWfsqqq6w+vwITec3TFXFVabRQ8GEG
06IvG0ISNUxLDNqcP0vFDfBA8LMVs8iPb5WsTv11aNVcZVT2J0eeIRciOA0wh+QNBSS1W4KRBo7c
D4yYWt7rvS2cGc8tOlDMwp4gDph4rIJlU5VdsL6V+sLGRUe6ALgpXJONJ0QNOlxR9bzTllbQ9mwx
NibAK9ZkNrUSBydREMOEy2XFbiUEjgX/yETktiN0QJvOJ+P0cnUSs9mBXPnsg21V2lNEMjde+Ixy
+/oO/F2dJhanRCPi9N5QfdxfH3raONSy9OvmQvHuLlVGxRhZ2vvjK0j2eZZr/AVMt+bgWjx0g8yO
riQJRqmS6prfC6sR/d0P9UAQVq1MpIuN0LfaGry2c4Xvczr3Kg/98xkyEvqhyB2Mvh0dujgV7UJ2
BT8oSJAxRSYxRb/X6YJsBEZKu9gy9B56m1J2g4sHtAD1afu3xkMgqDEuap3qIb3L/t+md2k+rjxd
FingR+zf1AxbzVZSuEXpA/5URP1B1OdLdNdrKo5SB4VgvfhmF/qsjZGaViAFtttYnflgPe4pm7o4
vg45E4wfrQ/+oKy7WSwKsayMrctoO8q/6nHVpPjGvfO2tM47XFq13tQzfGGXVzNRRG6s2U89QZUp
xNXPFqmADI61taurHOv5MQac61kjq31lKiCGsWRV43OkSmaLqFzsBkzMDPR70VQSF/ZA6vRUWNdO
w9U+K/hJ+18sVys8KQG+VUY5XJsOw9ApakgwrZaiJKpLh9ywe9WonDMQWx/bPaXqe1i/rOgmZvrh
Gavg/z5zvO0alKKwceP51ROudGB8E8hdCWECCuIHDPHDHWiL2i2gh28m5iqwd7ti9dp5B+g/S7+9
IL1OvT5bfSfQLE59VKX8TjRCrH5+LoleC73TWXtsi8VZaMADaLXsW/OZrurLW313G1yPXSg/o3DC
ifeyEx3BXyUsLmImDtOZvmO1NP9PuX6vJ7tfEQqsVoeXWmB9xkFmv1aTjJKHSUhc3qdKRVg7rkx2
BNL0C0k24Sgkv9YIUNYtWVNbVWXy+5E5p4H+hEGnQYXxojbb5W/YTzSO4RR7ZnT0vdxUFO8pBH+L
FSNl0m3zRWwBNQyS5Woaq/m31I96FZLKra58ZiCH+tf8/e7nJOYGAt1/XHbY+7m7/uMut3tDvbGj
8/sC6AvlBk6QlKrpyRebcBCWCzAIbyWa/fcMrq+BO6ZLAVteK0YnPu8YN3k4EMB/Ufk8JuRmccq2
1BtK4r5atkVrXKlzDwu5yJGEgGiEkEPpk9sXi9AmHVFqVFB0ScHv8V45FOWy2uDGfE127j/7PjxR
0Ds6KZ7RDfBFUT+FuiGWR84YhwC4OttHrcP0BfUcaIhDK7ecb6fgY1weTRYPlPvvoVfNcvlhUAwv
PTnMKMNGZg/dzYjrGVcwEZZ3TD6769Znl5WjrLc2TB5gixFwtY0FvlwsLO2IdSG218i+h6bg6tu6
3j+V4RYYS9QMCHCoph/xbpud5Fb7yRXgOY9IfvayssfyMVAHZbDrbQvGhAn3lDGy1vV+CYH1q/3o
JXuwY/c5wRELsXCMYZFlqiOI1qneBDBqPT75bRAvxMDskj3S1Qg1pFje9GXcf3GLM8/xHzX9kTSR
e7XHHwRKCwBVl4PXt3B4i/+n5vwknfLlEQm9+VYNymkca0nY/XzWVVqeF+Hz7lY8b5g9PeYRqHoH
BvMGFJKfY+Nk9NYaTv3EKrnhxk5223+a1rH3ue0LeK4CcQqvSKYB53JfPH9VHWgTV+PaWOYVh/Zm
z6YGHCL4JB7XQkaCHvY1m8SjLpRYunRGCZdFgmt+w6peQlxSDAJrFwdyRMu9EDObURBR0EpmjfbZ
55fTeF7wA7dP27k7gVVoJJwdpKj1KTiaOXhK/FSbUMPnO47pNB5Ui3AoqQdaoMJh/aDW5l4ijXKa
tdD9j6EvDBig0ExFSWilLZD34iOMR3cIWumcxBfGtCuTU8H5D42PJXe4EHoSlbWZPi6aw2QSuiDW
nqOsqKmdTbaC7+suf+aWsfixmswMonRzj7QOTAbmGqVXuD5CecDFWsKpas26ChTXp6kpM22z9ycU
AFSg8A68c1qoeWYneKH+lZyQxSIyiCD1JY7JgiXVa5jAI9LrxQnM2jR+y7F7Aeluj5OSDGplaNkE
709/qejo+oceqy3+RcUQSU14A7qDcsYfVispynsdTMbwoNYo3mclNC1VEvu2VMqPXSUUlyQMfib4
2ErK/DXLmkeCdB4jQ3OS2J/6VQEnBMAOw86H3ySfi6mxpRyLkbPlQofWvGtMfgB9VCSVvoCSdk2l
z6fbvM+bHHJsYirHPCIzX6js2StIQFsS/tCdDMbKW2ni4YdUwwB9ubQVMp0ziVmlD9qm7sLAiy8T
zA1B1e63uJRDNH5vi/2tw7/rgvWIKlzO59x7VFcf01Knp8dprLO6rLO+uRGcfELyrwA7yPhbK1tN
2oYLNIb5GlePLxsVnnDO21rr5MNqODCJyfvEWng/fhKsJJCkOkNPRaKn8kH6WlXMoeDTJ5sHqE4R
upIv6ZkhMh7V6QKsdM6G1XcdzG7MJJcZZXfjs1XysK8o8KLMCCM3ReNbDhrsS1a6557ZUdc9bAa9
CKvm9Y/7IUs2H67lT8FCKsRo2iJhfKyuoQ6OgmlayRLt9t4d5WP0nmWyYAtmhCtJkwun90SjVjWJ
ajvabCyw/3GLL7ZakAV4ftxdj1eWMx3wjy0vW5bArJG6hSD1g0W9rK3G9GM7Kx83QLpVeywbbBtT
Vymwi3WIHOa07A7LM14hl6MpD2R2/zadtvDvo7W+/EWQ19jDBKswdGQgGA5FZlmCmM7SnHi+4pxp
GnZbKK5tgKCAFf64egBon8nDuPQePVDQbdWSAHo/Yk6eJPsxOJdyeJd68524JPWpEUggjpCPuKrt
QOplyUUZqx9tstsaFUBSfhHGvuu9v/ysP3oTRAZtypQ6cOClO6+MuoAhk4ryLIADn8g0Hz7nNtlq
U+gQn1L9B+UnpiZz+KOEy1BEeojUpPcqmO6C+9Q+aVIGrYfFvG3u8PmqIVJ3d88LG5C+Y+NR35al
SDEvCdwzwv51ojp1t8CCYqpkGJ9gaZrKCKaHUhkN3M9j0zyQeevxtKhNMp+88IOL4DhnNMUStk2x
P4dBzi2Eu+EFNIRNTZcCK510Z/rtd7kQ/aKxuzWkdORy2Ymwd7ipSXBsNGk+LdvW/QunWQkaGdGT
I/gh8OBvdtx785BgvDDB7nUpCf1bpRI5l7rD6SnEXGTn4l6PkQ8jV+E3tcarwc7juPQiQKB4Zk9p
PYAw+vtPytR3Hs/qVW8mZ6AOr2AqPrMzUUBPDEZrHgfZW3OvzS4ul6VDvb4WzLdRbWGhcZjO9Eiv
fK4ryP4a1we7EWDMvDteio+RBv5IScWGYd4WzAknrPbb7JStMfh21jplsQzsW2vJ4Zvsryhd8PY2
Vbm4WxCItGz1vpc8JgNao8nCNeDdxeJ+Y66D4avj0rnDs+5C9K6VEpcgFLulCvNiCc5XliiJjGUW
c4WOyfedff09gDikKMVNX3a0wH52BvaN5TOUHlvHmyZ5Djwiah+HRgaSeJiLLL3Uyq1f0U09pbws
2cYeW2woJcmXBovEG+BiJxZ5afbUgW5hvj6yBM8Q4QaD5iKjH1plt4dVh3PBRZ8fPpcHoDg4Lyp3
dM2J5Q5qLyRgr9JYxK5NOh69XNJxSAz6CbQksGTnw7bzv1nOaKcywBUqNmlwJ/GQ2BBMyOmBkMpj
F/pePVm38KaDJe2EQKw0CC7GCbyolETFteibANLw0nWaNrua9G7odzK95Qr+UEDgpLJhxArM6WTI
Fm/aK9vgYT6PHcHmcG/iQSUZhfT1iGYA37pJAioFke3K7Iindy5PIbHQiM5u5te6HOBqliDrDTTh
2vXomkiSQZX5YBt2NsR64grqGS0jlQtbWxWXvaMpI8njjw++Jnkk1kUZD9CPphH4rwvpxcMOMBNh
HE/ifUYokp6ZzZYXq/Jauy1b9oWOry7mA2BooSCnnTuqVaQTJdD+8DckeZffQmlw4UF4MU4JcakR
eiyr5g28xfU/BhmJdxK2P87QdMFK7mDXebhJo9SuVIGSLEwXTRmPbNR8jgPpiZn4TvG+fggeWstc
042R9Su+Tm6mJAYhDgsuHyO3d09cOnU49SKDSqEWfMcrjWRshcaCgHFp9pwGvCjHSzjS5a3gsiWc
B5Fh+XflcUMNAPp+xZJC1P2Wj6vaZwz4Brm1v/JWD5hPTALgh1SQctzdUcmb69vyjhCUDg5EVyr0
/80qtk3HRTuWxJ6ZBjDFiJ3//ex1/8CPTSebmrSnIHz36+zFve0GdhR1SUn9fgiaBazzVwNlXGRz
StKEOu3Isc2+RHvB0f2udnCzx/NbdlDbciAh7OZ0scy1kzs2yIWvdryGXUBTB/wzHSASOgVpqGrk
D4YfTYEPaTkw/0A7qxoQcA0Yi/9HBx6AaXFQeU+d+/YwXnJiwHounVpbAkEfxen941T2vhLUAZ3R
ps6B1b082MtCJi79Apa8/n4Ph1VDlIdmvBCBucNN92sMMfIJd8FrrISBcPw7dHzkDeRr0FjiqqUf
uhGzr/69IQfzUc9xmBYvicNUEcoiPy5oVm1tBgPxJUPwlI3NEAYuvy57yAhYcGrNvEDD6YLowCPI
tfQ1JyVnCpKj2JczqV4cbRmFWj0BLsL4g0CkJqc/54Yei8W+LgK6mR7si0Ga8XbvHaSSFy6DuDt9
ZK66hw8ucKmCN3bVX3W1TWkRSkOLhITJ/u7AWQGrXiBzmCjHG4VI30wRHNfJ+XuNmjRq8rhGsQao
6w30XYsXcoAlAdXLYUrrly4s6ldwpVZwrUTz786rM5YaydVcX4jcYhBWrcz1t6Lkiu1ZBK1Ze86c
PDee3+vC2/6QvvmVDhgE9nKIUhyTROj4vOakdUVPUQRU2TVwCWhezwVTURDZkc9/wH4rUgUEqf9E
olfK7x/5eVxCdMbouByzf0SDPniRJTUTqpsc1AULb9eS2X7nkNDXwU+DbZEslbxWxm1sGTG+1TE6
QCH0KKqfMDRkYVo64GT6zQjc+n+06WuIkdEUpCi3lyZzTE5F3+faA5+wozG2uB8Ag7o9tRi3Wupj
oyhiNLdf3az0D+Tdw3fnuMpl0SeBbNNXGVx2iJIm7o3+dqCHwqBZ+2WP3RonMRXYK8V0zzotujmo
YsMEeJDvqJ/1T8OUdXg6dT/SmW+OoplM6wRM3IbAjy+v2r8yLHado3NZLnAhh2qkE2pIU7LfFsv5
SAWFKS0747UK278C4i9qsQ9qFdgeAuq3Z/7zaE0a8GzJnAfhnZkQMZnJAirbr/ltX+u0RJLagNZK
DTvWdtFPvOL55oWkhYtT2qeqTlm1HFT3/FZEBYDUoTSONuyrRmLAUMZCOk5fIuB9wjypLyeCtLkr
OjOoNJy4Y5uJd5AU0y3iSoDMW5Fz2LlfYSGQNFJTysnmCYvajbI6Q5QSI/wZqdctfsSTxOtP4Ghj
zRUPLWOK7ESyGVlC1epBNPv3ZCOwStKKZdB3hn3ImvANM03kwzgw8pHMyWgAK7l08zPgAOcvgk+d
/PYinJ+zV6r1hOBWtwD4lQZ8w23CwMx5NEwkCeY+YFLhaKRzVxRnd/FsaW2QxZd8jNK8ZkwQmyJW
2/duDGurO+J9mNLGI8/+hJTAlSq+1Jd/We1qT3sO82Md0kkxbVbl742PCJ7jmi53hJdttHeOs/xS
PfVkXWQpVCIw7koy1lOszsu00yahlM71B3iPIsOHno5o8LJYKCOLvKISI2ZRBFkNS/6TQc/sLpdL
nXSkYeyJfXrIyNaMv3KAHiFfIg4jT0HWYqkwDDmQSgjrV6teRmcYj9ISoUTGSl1dGAkx+WrBYBjL
R+L/8m7ASWfoXBoZjbZb6aLbv6NhuitGvPMRAZ6sIvEm+b2epSC5clbxc8UpLIG7ESCex0YqOT8Q
hgKZSkbsTKVDuyJlfzTDMaNLI92lGw/xXNQHaip+WeJEqLPevxu1yozeGOXyktr8GWXd58ylA+ez
7CiCy7SMzLq3/66HhO0v0l2tGe2orohJRBRL4DGeYX2zTltgYunk4QTp6pnU+15QaWHmdPcBottT
iCn6phrrC2/zl6D24W1JrLP5Db9hLQQey7MhQXfV3r19LFgtYPITzP3J2J4dF6GRcVJ9icJpWL1n
LE7URTr87l0tkRWOJDxtg2/jRw8OhhTKKl7T+J460wLOKiABm425cmGsIdWTsvA7xZgHfUGwVmoa
2HmTTP/RElwSmzOrYK+zATzGdNeSY5oC0gNa9l5mMKPagQHYiSjIL94NHrGLKHW3CYnXgXLU1vav
fKnbXFUx3NwSp6Imk3/JysCL63Egi5vG7YEj8hcgeCjg5xsKZDhSBjwMfv6lFwoU8oyeDU6FQtjw
1y2UIu9xtSouesbo8Polu5zfADq+is+ZpXkG3GtvHApAw4jxsFqWO/8dv2aAozyLhnsDZHFCoLza
IPzop7kHoJzgy1Sc4pwuH9qCm2Lz8eFfIO9fdr1xvuuYDaX+C4sBQcGveRM30e8psrBSzWws86JK
gRE7OoTZ47hqgpL0BGytAuicGaU1KaUTGrLjQUOwYigWpCroc36Mi63+oxESf1P8BPpOb0Aago6g
65JwfOCseITeBT74hkIxeUyR+1Lgu8Dkk1eiQhzBTVITON7e2GjZ2y6E0M1yNYdCPkXWY6HnOSRI
J3Lau3K/gdyfEeXrpauNZCF+zvOYzrbb/JHkacrESRJeA/GxNW9A3yIqMyNo3vKwtdxTamjgJn/E
NLScElInXVdfzS+crKM9id9xmn2zyZhaFBGxQFNCNqcMc01rI/Pe5Je3GmoDiGqMsTwbtTG6xlI2
T53ll9Oup+YZZJcx/cY+ihKODV57ZJAXIdnzz506ab6hm74ikvv+APkHHp11+zGdamDpCUm/KTDW
XbcuDtdXGFaL5n9ObJKtGA7r71nDiup0tI6K33y2/tgwjVBb+708ssvlzNr7fQAbzDW2Z2G4RRrz
U3VqSEEba3Y+97yz8M/Ox2bPhFp3UVcqkJI4UGezfFKsap3TiB6s423kB4Yz/dXV2TH3OULCmVCn
4eiBVoN9ftPg4xKDYWVj7B+TdnsvY35tY3+h1OuIgGaXpYcxNaXcKR9Pu1S3FXNiJtSjiCfmWN/x
eWdQm0HMG2/ozzqnjSOIm3IgwRGBmkMcWPbBF7DMQwidnb4ucwlH+80PGGfQHDikA8Z7y/I8zmp4
LgI7dSUV6u12Ty6ZT75ZVZEtqC5i8cBrk6+y2yzoxLBHZq7LF0+CXzNNvXQDZ01RkcT7mlfD9le4
dvXpNaGy71z+wuTp6U7NsPFP3uzHb9fzz336b/dNoUobnOHoetnm7VGhqssCu2HWhKbyKWcEevp8
S7RL/9TRqavpIB2L7lhiX8NPek6EwUcluO7pPtZ2ZlrcL5ZXUPjmRS6YVZCTKu9Gvwjx85pqyKFq
E4jDgcKtzxdoLU5bcYWI4SGW/HEKMV2vtLfnaWm5S9EOqB7vw7ltvE3xM3UeW7gIeXmy6dRXhoJU
LE5OnAdkteLOzGSWpHe71vuYHjmVD+5AkaM0OLc0qOK4uPZLsy+ORfE/amt1MZyr9fvDfmc4aRuS
QMRyfcva+3dKIP5HvQ7c2FzYslgO6mVJDNvDSFitbV4XyUNDlOlPspxScwLmtH0BIWfv8TwXDcTE
uM9iV0fOa/7qzEr5PEXPn4EFxnV0bxOBGm4wtPUB06Nd8qXYNhx5YZIEZonWd1dVf1i3mHH9Fwxg
DaAqboD0DoQS4eTw+cm271G5rSofoh7XTXLfkZrT37IGG+fTHi5m5PxvZDGg+i7/DOaUGjb98967
jv7pBI+D4Cxw7vN/IyJm+Y80nwG7UvaR/0k1mHOMSQz48STNziqXWwgmRJXDFJz5zWzf8DtDGJoZ
Pegz2J+KBOnuqAkZPq3rvgjqJl0VTur8Z0ryEruNTT6UoG3y1b3DUJjtAlMb3F45L4QXNWyfP8gg
s5P5N1n6k/g1dSGIARnqBPaTBfLwm4hkFSR3jx+sisQ/70Ph9dgD2rrz37bsIofQJpF1E9DIuNah
a+9uxhpBsFiWsJzfU+hlDKgKRBexlmemGkCf7euoRrxw89OxjHCoNZQI6ANTonRmRqTYGl3MTFEL
5Lkj/ifLq56aha3RvOhd63DyaU+G7WfDLgJaOSoRlT93Hq7BFUA11H9CutWe5aZoOWTZw4WDw/qu
srVvav5AleqSooJDiLMz3oEepRuAu06QmYmAFLZoZbrb/rWQkdGaSKMym2p0vXo2glfmKZrO+opU
6a+5SI0bCJtg0lvehsNoH1YfKhPi0cQzw2zHj7s8DrrBjKBfoRqwAmACYaBgn0gRE149r8eexl3g
tlVk+4YRID2R5yeFh9JtQXxDKcoL9gDJ1j5pivwyU5R+uZuEUf5qpzbhw0oeGkm7Qs817KgENxcP
jRYq4rjrZ8rJ0kF49gBLFyLp4VjJJB5JJJNL6cbdwu+u+nSiLdL4FL6PCV7JrggTMlqNQfecz3ZB
IDkE+OTp8r6B39Bjrn5k2BwPxH0/71DJ0ACajxD9so6mTOw2cTRYVhGpx9VJqJTownd+t+wKyKJg
h281KYQ1e8qQrUye6gzQxfbi9crif+AOIGqAf186IExzRCRpKC1VLczwAQK4++OPI9dNBuytdzcv
LoU8z/ELTkI4mx5Km4wOCdVXWnGnc187wmLhSk5ioTR3Sdulzee9Qj/Tl6Hlww/cr0ZH34VH9H0z
Z7CKdiagphvmr7raGwRhyu9+AYdEAAsvU12oie4jUJ/Uo6AFIZcEnO1dT5efhvk2AyQUoKB00Ri5
E4pxPkiSpYmJu7QPgmijRE3frxAB9yVSTmEEbnOn0S55feQrWqSoqLYbG8d14HVQAp1f39zTui2y
da82MKEZLc9pfPQ/6lH34KiKxLhjcx7A8iJZmQRsKgYIfiV71Eo6Qnp5i8/eV+qDP2s/+2P93N5L
jBuc799ZsWDdwJTDppDre8LGLrOfWIjGmbYza4EMdKMpy930zDWfQtI3dkJqmfxdKOguKZQeRBfS
FLcgL06no5rMboLXrTvY7F5STLtSzl81yvnwhan199X9RwCWQqWkjXwQnAQut1kAUQj0ng2Yge6H
kmGV7Sp2EhUWCL1ha82g/AiK9m9gJbthLu4kKzgMUFdqT+l87a2QPXfmmihNUUWdtqBjg2KwWhg0
+uUn/60tGuzy7bWZAihSiCnums00IVRNVR+9RBY3C6QNdEdIWal8rWCRpfvVSge9kB7yBqQ1N9ID
oApVwTPiTskYQYpwJSuro9lZfY8UEE0iwfOXG6wAIuh8GFPrKOztP4z5Wzx9nG27Yk8OhhtdTZxY
U87de7eq8KU6BwDgQnyBthQrHkajYZ317UfJ2whrFMfRsYLwoB4EAjq1f8p8Qvym5Qx60m53N63j
l8JUMxSfO7y1Q/mA9+JloRkXSqfAWrZgyCmQZO3dGhSAsdHU28JZOFrMII1EQNKLMv70rmLPIWK+
aWTN10cvoq3EwozyiSUBvv4++Jqd6eUt3+Wz0TGOQjFR2S/N+vWq/ydgCb6bH1nbBG4X4jEbVOCz
QQ47Hjp48I9gxqGGyLD+T51yO71w9MDq3/kxIqaQeIZxseSkdV28XnwJjpzy+LaX6L/Nqal530Yv
UADzwBKVVAKwu6YUqx1JCHUlpkkVFsN2STL1j6gSjxK/sF9K3US6st9VnyfYHJ/wlQIo+au36cBb
kos7iqkyp8F5AJ9OBVq5pQte2+nIKJjHQE4upjChMIaA4o9KgP1/rrEw3Zvh8LT8BelsXx6zjX5R
IVT4TDcpywa5ufuYL0iLRmTEJuzhA7GfZVLIJuo6u3BzzqUguVlBtBzlRhDO2rPStO1gM+N4EDkc
ZPcV37Wl5snAQCa7k7T/91RVoMdlcLcS+G3il9v6+kd3KAfxBEGr71F0twEBhdEXVznhmtKlDPvm
G3soqWrHzvzovJJiLWIxAsPvsFPtm58oJyui9igzEn2HXayHkUpDiOpYkGNGpQ6fGvrOVeJp7b7C
dqf9tJzqG/xgpCrsC+vwRZFMK7gU2yjyHLVOj0rouq+X6X00J6Ea5DFVQiI2678QLNBvmB9Kb1Wq
6Z0WFtXSbYoGogO2H6AebQIqqdwd9fVt1cXkE9XAITdPwBH2a28VkgZ0lfr28OcTUDd0y1HXtx+K
OaPkmWMdHCQIOH1/RAovsnjwxNhqPTJnXK68GsVBsZ21aIGfzlvP7mmeleUGKnTylKvq8EbgJq4w
4LSZpnTGj9UJ41QrsJqhF2yJqGxgK24ckOcGB7nhmG6Fisxk7SuRJ2ZA1UkYLPjHM6lP2h6HV7eO
QEs6Ssx4kZCsrn4Erqa05f7swtxAnFpcx/mrYiaTbK6KMYRKvjPTwkLfHkowSu79/iQ94BU600tr
E/qj/GMXen6MvcrsWqCI8mYnjyIWFGzyQqX7SGpwOZwy/cDzhKL3RHJKzZnqZokkHX0NtzlVTnNH
B5Q3o3ro8grGG2H76oJS2Lez9CNC0hc1ahwEdFz/0Eygv9T3Ct8ih4o9bugOnhCAH56m88JTu2os
HcbFDzo/4Ys5gR6xffOThgPsFo4qTQn5e49EWgpIWNY6B7zd58TbCMK2DffI7yRwy7wZ447cbh5f
zk3oKoPwiVOPSB8wPRjB2M1XfoqmpOgZSxYeX0+MtxP27iomf2nFrDAsj8eq5K6zWQ+7uxzbzzq6
JgNjiA+hc44A+49VWmVCBCA0JiRO7pYt+HtE7XMQcP3sGheZazhQ37n0eidwA2DSsSSWPLFTvoZl
ViIknIjeIvBoO0ylQ3RhtnHp1/dvAdQgrMzdpPXs28mC6QHzSYwFTXhBVGbERjWx2RF3DCt8JyMc
oR+CTg+Y600077NL98YsZD+iQlw0sU90u8W5sNB0iDSFr62lYeg5Ugeotphi7JRXXHz0YcR8zupE
nUzOo5cSyzZlwXELhIZWbeElWsAg+sPo2MdBXiIk4oLwMYcsdhLV2YdIUXs3j+5SIQH9W8+g3ZGn
GSdK6/NA5hRdUrBirmFJKVbnPDBXViRP37Sg+5q2D4rVINi4cRRjMSUoAec3XASeXAPMKOrzZcSo
eHXYtPfHGZtglBPn5kY1A7492LL+FEBdLv8of5ZqzCF9j6bi1B49WWWEgcIT1W9/X1F9C9JfNWpk
zxwHnVJLLcBX+l5I739s7LSIiZxt2CTW3Fsi6iMmx4OLDkCMR2RI7Y35Od69o4JOkVPxbPOxxsH8
jsnlyxtAvnp3nFDGxt5XWiyJJBksCKxLUqD1w70JCu3vNgKybftldvps7bYKE8TntY8rnA20VUcC
06GCxi874DpOh4sEOeOA+SdzltpuTn8uwXIHygxoolMiN8r0FQyDGoOlcmU19Ubct/Plbvk/XGBi
ebuJYlsvllXDoiNlEl5h2eXUMTztIQP0wtRJKMiCzqS4WhmpfO6l3rst5F2Nk/Nj9Ui5oSrtu9A7
6QdRq5SpCLqMUTXx1qZLGTwTKm3BY1Cbjf7smhxHVXaNLcU+olkYlP/qHHmtGZ/b0/iZ7uGgT8Vz
r8O5YCRcrN74xE/u6BrrKXVI3b26LdfegwP5kDPC4jn/dq4m66t6fC1EHB36nF5iA0swu73c6PRV
11MgCFXlx5IG8MnlNKw3uTI74n5Uuw8zGi4kieFjfwJ5IX0r0GR8Hdd8wI3Pslfs8Xcdy7mTL7rc
0ft0DmhN0LXEN5qXldk5+A8xMVTKBAHZKtdMNuJev9V/s5zDWaJa8S22HHgKl8UWv8r1LPGH9Yoq
qsZXYZxyckJpRDtr8OoPz6Kur7hX5pwNk0vClt8fsVwelIZ4X3UbiZclI+e5Vh8q60L7kqZN24WO
MqeIHCIkDNyvJ7EfWMb2Y18eJjJXsNIalebKl0eZkBeiWxml9WciFnsOwPgmVrKFZdhDflDUSLZe
DbcgpGPhpDKUhZ3CgCM7d1ogqd8ij/CrzFULtpR7qA9tc7aJkwLPKo/i+FARpA3TBPXZ4zjO5wVM
QoszM1aVRoVboHlYrCVgk6zDkQeDNmwAOleShzvKNG326O9JHTbDx6FpvgS+vtZGeNsB+vXw1yai
AhKpg1Rebp1UUicLwDGOp/+dHqF/yrUa8snCGVF5TxQAddUZBzH7x/09jd4c8XXOCnQQAtfD2YqR
aJRLEnQbdFzW7ltrSPdDUnzkgi7NM1yCTtnailz3/PikwW6X10aofKIIkqpJgKOZz7faGqrAYZAi
eZeJq+coi/eNL53n0yJY5QHVniTym0yiLtxvufZE5g38prtE8VixTIor4YzGWHw7YSjQx2IQpIc0
/aKtDjYQe7hG1F9gkZNTcy0tk+wcyLrfL9ywUKiYxEsRvpEqcD4QCHQevmQ1PmLd2tWJBCg1lwif
0AjjRwsNx68mnOWRfc3m0rBmXp8VBtUfpC1aNmGRVXHp7OWf5D1h5oBPlegYxZFOclZ/yYTLDcCu
FV9QKPVA5uoDP+MtviTex57XpYzJ7EGnWWaZaxBVbcN9mHea51FKBfVzoUlL8zgoL992OiB5Xzbj
tM9Vk8S+4KjCvw1RC4MvyieIjCmzCsex1Zohwk44xO2Sr22hTo8JwfEQIokBX97BMidAj8jWAakr
ldBlTlPddC8EHjHetp12DnXKnAVpF4K5sp3r+x9Ok+v7RkeyWBw8y5DRNlnoTTZCJkROpPr9gk/M
vGnAhTIzgVeb8atJIHMP+Mz2G2soT32b9TXq9v/oQuJQYqDk+dT9yIO/eSj1D3sVJcm+za8YyRLl
8rf0HMDGSdu5NoaeCs5/mKkbLlHRRBmpE0+953mYydl6a0LqdCfYrkU0EndUSDaZm0eSKkRvN5aL
2zTCwTfUHHEnvdSqa+Q26h2b7FJsUzRlitcO6W5bUSr7oewTaJ080cZSNEQJjHZbwVmLE/Ayynzv
YaKWaYWkLjH7EKtq5dZprv3s05laPu1xpsuwFV0APYo37lSKN8H8YmLf9fT2ujVOEXl5c++zJQIE
MAPv3RF+EFecX7umGdWIm1llt58ShjMgKpbboVCDDhGvHj4mYBRNDuEpYO0zxPSdtYmy+tiIeIUU
NnaULQ2uRgnpy08qLbFxATyV5k4x2he9eb/glDwyjyfXc7BhDwTWyP1oSmuZ1+Wxa/xAlEcddqKv
tVXktPxqk3nMJwIGt2DzbsjEyfq49+DLt1yyQp7wMvTW+E9D3avTKv26HEeABElK5LI1zVXjKt18
h3ChH+bp3cC6mcqQr+dWHFe+GmywRm2ZWT4aUrK9p6a49TI/Aql9PmTVTH8OA2S3BlPQzw1c+jxd
AjrYMe13MN5aGfX2tVKi8nlpuV3PyfjizNrnY50qLwF8FsZjZ1yRrlvZBCG5/V/qcZ/E5E8ZXjyN
NYq4vVa60Wc8d+luQqEehZaAq2lG+twNLXTqQnycycT/sfTjO2z6ta2essSdn68L7sX4fOEshY6+
vQkbWt/51im+oPnHkPPc+O2BLFsBP0knI65RhCEB2dtF7sWjneqWsk+DCSS7TI9oTOFigUFEvGnl
IKkb3qXVf0qOevusiQeIHqj5vJMuZL/R2ijB8jdbZV6vIQHDilg4hGQ6G7ymOFF0g3Kx87MnAPy4
0099ThCXRXzXrZ/p2icyBJuKIRIi1mRIrsAOPDfGHOBW6ifavCW0++UvPdWSfb/0ytQq8k9fLmSQ
5rRZHSAdLGbj8AZPWAOCLyjWSUMSuIKl/yzWOnCXnm6fUvaalflDSzHmjeuz1fgMTgfz82YSlxqU
x9ut/YRcoHuaqjAP7N+w/FUj+8pi5Eq88sEqy1tVTmVmPOr/dIm156IlO32QZmKShXdbVfOxMYVS
AhL/Mc2F06NMTuDhEJPr46IiPG6uom8p+DV5HkDyV1XvNgD1CUrnpgUZt78mV4FrUamhcMPz7LpN
HoNd/HyX4rN0nG867AmVnz6F90u3QdwTeT1Z+s9tXGhuU4t/Eufk4/te6jFa/Obp7Q07XOQpOMsS
9A3EoipCV/Acy8fp2Yf84EyXgwXITACciad54QQKsFQJcwr2pwa5p1p7lqJnrBPtegAkq8jncw+m
tJlxlp+lSpRwsetGe4oKGQZnEFbjLQ4s9TaiaiIytLY0QROL+nT8hZevoPvXldk0H71lQAj0/nu7
QWsQRXIfECxBUIYv1Oc0D6lVkdtqWLZ6Wr8Clyk0Q7WbXhiVV6vbdmOXaL0EfecasDQ4uOoqlwN1
d4cDPUSUIFpIEPWAp5KTGFb7CVQFsJ/SXREwURVD6LV8LsYlL0NOSlKkXCR/7CjG77jQq1x/ebdu
64NajuqAUIARL8SQ8LmH5eD9jwW1V5EoOmuPuYCnMbNUzvuHytHBAF7yMLnvqJKlKUB/2VsqP0Eh
TB/t1MwTIJOTutPK6epfSmfu0NxqKmPDoMZjmtAr575RMr5Cwp2UFB6YJx8FyH22MXpfHs631Dt9
Pjy9Lk3D46sblzkBG0C3Nv6L+YGmPAHtMCbl76hSNlS9o27qrV1wYjhYhYf+lopkBPM0NRwR1SNh
hlHx18ZIDShgMm8YMkzVGTTx8snN+XG49nauEVlj0358dhVPP7WHvPiBs4v9L9nZC1XzxVX09NNP
bYuCsEi2IK9AfEU6oHeZoAE2ScJQMRrMekGcTwTjxiMgQD0eO9UNBpQUqD2OJUy8WX+Hru7DQlvn
C30NyHrg8bd/ijWfqr+hz/zeCPetcHZelNe8+fNmZmGSiJZAhncg8E6Pf9XMuin68wFbDEu/YAVQ
yfLFUSl/+gfSazmykX+QZvSs994geFR2OU9bRsoRRN9S8hWy870YSar+tA3Nxt/4odSnA9qBD6XF
IFYm4oPYTcskTYqFaHHo897uISUafx/wQRHOzzjIp3wpPw9Zq/lIzGNwzUJnK7NrRpjtWQiu7BZv
jysSpZOPwPicwCxKmNWf3vUiTtX4O4o0ZnqrMVUZhstwXjwrm5AGifSttABohiRjiHnsJ6kgbs4Q
z2V0VGlXdnUnecyGaCnYU1H1mKvX+IjER0AgHNbMU+i23/qRRpTLDSVWjcVzHdQSnZ9kqVnf5any
EnMmq7YzT6MyGHNeNPp7/iuRFi+Fd9XuDFOd85W+OXcg6o+UdHUh6UkEx+dFvG9Qsk1bQyhF4stt
cFd/j5/6Au1dHtXGgvYtOY6HaFhOsNxBu1+c+n3y5KbyTHH4dCCv0YELnexGqeXEKJdKDhG6G89B
A3klJAi0N9FmovKjd1h7icQo8swJ8ZuaBvLAb01iTIz+KxSmcY3i8go0IMchtPnkQZwVT1jLmESf
JiTBzRsiktnSRGIuZzTXGa3+d1pzcZPiZ2UVxGzAFMkypy7kNp4Dv9kdRhWjuTpOhPszUul3+L8H
Xq1YHOSujIGqU+MgVokjvOrfjBk6G3M0DOMvKlgAEMEW3ValG4rWanLNczXgallryoOYb7K+zDAp
0HOSuMl6avff4NAIgDZkTB1JlROTeDfMW7AIgbgzuejbndQpKGj7caPuzUvyUgBwyVeBBhVu7k3Z
9azjFqXIgQgsBZzjFIiMPZC3mXCGYPjtsMGtibFImIsyXNr/1DlQied74sCy1SclDX42W6j1eVDI
Hnk2Ri/Jkga+yTupoZ+2V4fHc/eCCnDpE5KGc62oQzTv4qkW/9VqFzw5FiTsS/NLrel4K4ZQ+Ib3
q1W3hJvlqnHXG20uoLYqgIHGmYAqLIQ4nSj5gk8lzeI2S5FhXXgwcYelKfVJF+gBR9RyRQklDkYV
9EmbNjq0QaBzSIUdRdTjOIkSqbeqY7YpUT2VJn5clzJLATlEobY9v5duWk7RIiq4EceyjMZX0nJn
knYoTfK7ru8vUBU80okVvwQGZ1eQs7E7tXvLrQWlCfom/GZaPzQwLdhYDmUshr4awSz+seEg7GFn
Iz5/zGfA+cJxbd7RmVz3hIHFN1fZc7Z+9wyrO79VH3iiTYqqCzkb4B8R/FKe/xiBYyF81nO0N74K
nFE4d1PVMc7Y+YkNfKCPfiXks4shAzpwaS5OEionm0prMDhLki5JSu657f1KpYrmFBjjzmC4k+k/
5ygZ41IQr9mA5lD0DbKS6Y37aTQqwU5t56/Hgq+51QrcnkDCfkuaUlwajsvrGtbLWJNBJcULyn+H
G+mprQeAwDomEImQ6O1fllQD5Mn2LNURra3/DxEDIL1j5WaB5uBADQ9mbmoIXFeVq1dfKpLG+VlQ
DhSmZ2mwQfYja1Y/cB4+UtYh1fqYoJ72DMEHu9J6RyjntQXpYXZdK7hCFUH9N6+XYrG8uqiwT8Ea
ouf1SNsZks/Q5FRPgYcmIctoQCwUrN4PT51yD7BDcTxj13bVgeA09a7CVKRRoLeIzoeJuLeTeCzW
c2S3IeCDvABqjucCZrvi3CtJjq21znLYAduMQrXeBvGqH5KugMHE8ou3XST5aL4qBROC24g8ubDm
385iEd/2BJXJ10kbjkut3Wvzm+CSM7nSgcuFowAjBC8AB35pxeN2zde3hbCrMkm0R9El4RJKStI6
iQL5Y4eWKp3UA0aWjAurpWWqwxzFUIvpsZxw5hRLT5TufEqkyEEyOgyz5CVk52tdUXk0FrGMj9vG
QvAGPNnX4nRughUB1KL3mlDgecYh2ZZUHwuPM8G8/Y9ov11AfxD8BLh5IVOcuFOaM5t3I/Kz80z7
YqnS08+/gSBjaT5InLKsHaAVO9BNb6O0HDJ6MrxUepcyigJ44AB1nI5hKtpv/eILQ5mWmXvea+1B
tqxmjGsmP5oI0VuBKXCfZAWKSgA7NHWLJUruOiM34JUwm47QnEPS2TwTxIx1BuwWeJ6ZlM6JzEPe
sptiv9Ip1pJe4seHKvku2EIYSpMmYBZyLIgkrBCFh0G/RGPy3YaRSJAcKd0D5wHGpAd3fbdf7+VK
hBpNn6r/bHJCx7W5j1gQ5yQVC53IYBVU0Tw4uKdOklnaSVsCPf8I2wdG5PnkC77t9q8Lj0SDx3Rw
NsX4Mu8p+t9L6eA1RA0Ly3w83Z6bCFZKNpgFnjFypTx694UIacugr4dmwPCjnuC9zxA0UKhtM6B1
M6bZfZhsO5QuR/fTU0jnrIjbOg7fCwuFX5jxMsFGYFi880ghuucuIflBoPNPUisqFaC+AGc39paV
jSoq4JTu1H1uH2zcEGNeUnE4CxOKvP8RaVrCTdwv1nfj/5+wxiSmuPX4ap/miItrES7S844BRaqe
w6KUmPerGodi3nowBLdiSBFdFf7GigwbVhumi6knCEOtuINdFmU4Ylkr0I/2fPKU3Bpxx8AfKTXd
TWL6kIyp4NKw5FikAMrJxkE6IIiggPOCVX6mBrYKoJEa/wovj9QPc28UpFZR9R+YaCd6WbN4EEdk
SgE1KvBK2K/cAWNp4PE4GRsKiGbp1lCbj2jhZE7KFvSe1BmWUZrLp50ZCdaYzTEu1Y01dfnrnngL
kmS9a4+hqyYvmRQWkkWjWuIXIfIelkzo3/ZT8HTHvWYcfTFdJq3GGqjEc8dDFrT1oMbQDTkSwZ4L
XQlfALBkm4fpZrAIMW0fpwrIRWRPuu83kYpzxDtx5xrg8YqsN7XRdnHc1MjNXo3mv+fhllGaoyum
OhNqAp3pmk3xf1TIw5OpBDfgPm7B0B1uB/Oi7YE2GqDtrV/uHta1dsOLXZfot4dIkDVf5wMfkubO
yvzyZ+k70VwUsxaVt2bM8M3jYwSsJCRqDtpy2+yz9mTsQlbpj6QX7iYgH+Y3tHvdQ+DLzlt2fbkp
JqvpwY/aM+7RSynkMCmBP9e/KLrbDVr74+OTBuIFs+adrC9FrvzmAT0uW9JLR03XxtylcBq0yDeq
NhYIXGXT2mksAMPKNcsIkhg6sUZAHso1wyUlMazD8wgcnTRpLP7Gz6IhZtOc2NHG0NfuFImhuw57
1FLQRRGYxKV+9ummYrFzt3K6AOrxT6p3snSjv6xlbJ+kxsvGaCvpc3k3RFL1FZ1T/HX5Zx6GaBBi
u2g63heR4VoEf170kYYD9ZNQ4kDIHqMm7X3ipI8cYVmB9rzKsb5XVtPEmYaBzc7+3QnIL/qhptT7
RCQXcIrcW/GMuggySfRizRwW+xTe2D1r2qB4Nr4F3r4m2+UHNTz1Q0Y70ZkpR6g91WwRo10tubFt
7k0qQM4rRQOZU4V2h3Uf88s5wnbfvJmwoyzG/5jIPT7p5e1QeOQH+w7rCasiWwZEIq1Cvwx9LVsK
jr+07Eu67klc0MJjmW12czcP0ctotEuHlDE9xRuy2uMRfY/tVPcrJp87uUN7joMLx/QeyK5ZU0/U
e9t+j4MllheklOijrfJQtpu/xFHvMgQglx+HB2Fg3smuNpORAv/eUH/XNJfPi2YA5SKgIDk9COql
jtYy0rt9rs1rwOoOqcsSzUmtS4Qjv5dkC+yfw/7Hd8LxnIyL6QWWHLX9HWfiEqCR6ZHA7po4e/C7
PkzPQcM4XPrc7qa9VmEciCfRGjQb6ZSYI9V+NHQBtd+4xHATCc+KeocGHpjq7gre4S4k2B55fbLE
+j16h0lx/8bWkA4UXeQQX6/HaYBPcQ/uFkQMRJQ/MRt3OggbYhvdpggQnAznlNHMVoEBfNTZAZAG
db0/+FhcoDrDFiH4UdN4Ki1aSyQ7nFxjZUmCuqM+KPMFgtxUbUFFJFjAoa5OjzYC/iCQqxAqEtzj
6vDhUKiQ+sF39D0FuXLup6ZQqD4qO0BobJm+aLRLE7VytumTcjQaF9pPB40sJ0h422+DzaDLNGKP
sbWrwyk7wMecZulS+Q7BwGorLsPx/3dDNmJ7dWBzfZXxO3O4K8iJ4/DvkL5qEhCA9ty92NH5vK7I
9tE/6G03Ds57/1lbuvtRfucamKvfnDFZ4AJ8xxJmMgkQ1s0Tr1RNyBiXLYEsXm0iC1ZsVZHiOhdC
CYuKAQ+cwxWUc9NLKMiEGiQWE55u7Tv0PP97tQ90IfA4+TN5KeUfuRk1+UwjzzdjLTSfcs6rXi/8
KK5Xf3645gkJdwNiyVDbFVVpB0JsbWiEyTPyP352pu4bynFh6jrRehgz/6k3mI5ziWvdcBYV7Pks
1i/cWGqnGiQqu7gmvHRIQLuvj4kd1wGO9vy/Fse/6+9sX5ZrhT18mYS07TII9WJjZWysdLvqPTZc
+d9MJ3JwwHiB4HYplkC9JYpvZ5pHXb8YZkL1WcQ4uCUp5MFNV+XnqWFWEzeV3TZajAm9qZroMvtk
lTT9P/+WY/Ae8xoN/tJ8aeaXchUQ7Jo5cUL1tKMoLE67T4Id+Ce6ZmZ+gM8NydL7lkyXJgPHmQU9
ys3eK43TV6QZUZ6RlQfeoS4iNl8sjTpY0tUbBDFW1XHXZRvt5knsPs1L+6inub3jm3oa0wi/p0LR
vfWuaye4it1LifQTYPlYHQBD0R/81do/rMQoQNt3m7k7yY7GFjFO2eKybsRtRLW26LZC2ivT3PQc
BwAWGK9UHix9GeYrbIKvKIMEG/iU5/V8PLiDwvBPeel3Qbrusv7nwuR/qTSmOCiISrbHOnHVyiFT
amz4p7wljs5+DaBRmFNEbHNaPJYK7MFoKyPbBUwhiwexbnHiN9Gb1StRYd7TMB3vvtCmsSja3sb/
LlAPnkegn+OY0D3i04IXE8qr5o3Ul5mQUjA1tMIJ3yFofbBNgFhut4+HAjQnQVLTlR7Ce3PsqGBR
08qAndJTkuaPqd6z3K3xWJ/ZJsSJDY6wa4ZJh0Xu9alRkfijm8gPVvcEapPFSxZtIz17/kgEqd3x
xZWUhY8oi4CfVphv4EnXkis19c0geohftNOzWLGVxH7uLqtMpok0gktezIewGt6kNvzwtoZbxflm
M7Xo3WzlcZFgVYwOUU/t2xmwwgEGmLB2FRBRqfE/qPfGhwb8emwQ06ppxWa++haRjBtXQS30Afkh
/yYF15mqr+o2eI2p8E2N7RhYkF4XwtSB/mX53IXlGSAI44uW6ne+fYn6+A8p1xRX9GzRZRDyVw3P
HuJTeBX67Ro5ZXld/wpXq7olo9k6qbO7NjLOotq0JpHZ1Z7vyjdw38/cxUx6ZF3shdKGVlkQz9tz
NZ2epf86BCFJ19yiaBx7gk/JFkWeD+74vyzAOKsF0WffCx1Uo4G8Qh3AZTOxFr86dC9Z55HVjaOt
tb6MiArxZzXcQ4axGbAoLWf+zdUiDZBLX5Lserx9X5ASG2BLm4DnM/f1r+NvwRVzc5B0gStIXDJ2
hS5IO8XmBNgYxsdx/BU6B9TSDIAm8ZX1ZQPRM9P/M5Ul3ThnLJLlcSD549bYaOeZriGGtsqN3ITd
XfIXwK/yvY1KYRe9TgasYUPKLX6MHMrv6HGRK+xaPeOa0jJk2vv+7e/5+AcygLoJefhR/xOS5Eup
fkfuQyUMCXuc0WnYmj5Q0dEQGmepefIooNJQ40JCNUBbQRGfp/w7hkIOVTr7JDfuFZILonNprZ+j
DEk+nikl2bYcn/P4cVY0qHbUJqdexoc26cH4Weq9h2sEx/5WE9yWpGZZBAKpmTaky20flDSzQiJr
f/gRS8HoRR1UMOgaJMQ5vK18JzQnq96R+kIGBTFBTijBpfmXeS0nEPtfjkOW4tmogmkkC2QGHib6
t8Uyn/vopsh2iLdgqngo6EJTxVYLfzokS2XqodAWjtiY8sKKLYcJCZPAL/et/GmJI2IsJAor1J0W
hVIWiCLOBcV3zVoebuTJ3DUaQ5xVU1Nndi9P4PCc8e5qTXAQrP87UgXBWoDIxZ4pH8qiPlv7VIKG
NZ3oQrQYC1lCQSlFs3koCcXDuzGEc/OCTRAOZ9k/Ve4MOr7NgVUSFH/5dDvzenKH8+omHVHvn+f2
9oh8F7nxP1cQnrlL9Zozp7rPD5rVNZtME7jKyMSWb/xa+WSJj7ZystPj1xeTGWRHnCQXGnJVovl/
UE1MRGntdIxYc+ybKw6hRkmaywfnyi0FLGedmyamCem/v+Gvu0uFPGAcYEysQ+drjKofUZSeIJrd
WgH3mfT98WeAxjyz/+nzLc91eUeybA1dxcNrN1liRoI3slI4BMiRjoV2BtyD7yTuRZUt1KAgnzHL
kzMuw8Tgjgt+exLY3jav8LsP9eJPoThWh1dEAlTx98FJvmMKVprsW+hhfmnlKgFiZ5CxxzkvzD1O
Axe+4tvUPTS1gVNshYmOjdPimzZnMaycH9wZ4anhb/ZFec422XK76TXKeU7btkeryPIgecrO5CDO
ckqGCTyF8ZHmzhuaA3CaMcOkLtKJRUajRc3KbKNKNm62Y7dFzX4Xe/ga3YDgTA4UmgJKtR+jx8PU
uRSMHnrWVa4Z4V+1SLfybZGeZeo+g4u29vk6oLk09H9+g6mFwzfh0xNKLHmJry5lA7s9bbfh4nv5
n2lp0TzhftyETMPey0wtck+aBeTkE1HnFIs1MfnK7B5SekjrsGwq22befq26Zhn9hbxtKiAL3ahW
wXW16nKug/vda8cKIB5G55LLNDCVwMXDYUcN/g/axf8br1po/5gmBcWu1cVlzDesBkywO0HJ4uFK
1A7jiDkmJPDHQ1lJM5fqIP0L09h2QF2FXErgsFpaTTi4gFS3FXRJopCNWKHt4YQgRiyiF+CjqOkg
ST29yUtP2gsAACbcVdQcUBzc8+5uk1MAiZtYZozp09rIBJLb3VWMkes8XdNCV5Q6Htzj5hYxEL4r
MB24joDH+d8diAu0XaNweN1C/FZuwwsAWGWWV0WcONax1OYDlxOG4I/nfmURTtJw+tg9hxJ3EpVH
g9lf7CYH9Ph8QUBEnKsYKN1BLwVLkdLIzfciB9BGr36EXXJ+CQQjVg5YBQPEpiT8QmkHYCQOcsHa
MTE7BBEf41la8tIt9ZwUBxJEo6KwiqbU6zlsK6B5CZmU9HL7LRrz8FGj5Tv6w2N8SjZ4WkXThUeo
zdeeKBaJLT65ahgfPexs/6eAVQQ5GPlSCgVpwKCXXL4WHgNj3W1YyjkreXknNMyGAq3pdiZ9e+KE
6NTLyeurY6Tfcqq+x2s1riqLCJdN7U9JLJqlLizWwu1FmJK1Mi/vOvLckcMrprn011NbI8BQ4lGq
fVyWCWMAN2xL9h3Cqov26Q7nVDuGAGQannqHsENFkdCL66OlYek5AbmF8c9GIo0cKZ15SMaOimxa
+7SAxik+pa+X0HeHUgt/4oq9nYfAhIQnnOT0z8qiPHl1MLfOEqPC4AN445pgXanTwBFaW0GtY3RI
Dt21irYwycFqzia820y9OYj1p7rck00at5P5XN50m+DdGWHPIqnwPdMx68jMSDh0b2CftNgmd4ap
LY56C5yZrbbNiXPLJZoXz5ie05VQvNSw+UDXo/zFkF7HGKov3CCW+ELS6A1BA2ISgFhroHtZEjNA
UQNxoI89sl7d6gF5NIYozcAtAFzGTQFaSq+CDGiyNjRH1zOFXkqRb3qg6l0Ig5Gbkyfoay1dPkiS
Gt/HknfhrdtpSE7PYmMex4gGMu0tbmBWvq40gaGAjwU5iNNldC0nv/k2uzksWPm6KXw/yt0biPIC
THcO8Tikse0jpDUT7YmdeEubh4yaI/WKtpY6FexqoeN44ivPKctrLC4WfQ/KIlJPnNTDK15XKZGf
OI40O3tmihLCfFAJQDQ4f96nj2gXqeTGMsmMWR3od6/S9rkXEyfzzCul2S48rbFsjqLXkhcTkWXB
KhhGkVMZhhbJKqBB34BBNQBHNo7UpUtszARS/tgSx8D0WXpoCUuLwSJXwdHRmQiaOuy9p+LNbkAj
J6goPiaNGKDfguUHk0otd+SBYn2IoicX0FKCYgVTW0miDRF/XnnOqfg2LSZ7w5Y2XKfKkng1elln
JGuQIP0NIZTdkt31V2j8ndTKYFPiKEbxvTp/d0uKvU1+CCXIjDAtgzacjhwLphCsErsOUvrXwkri
ds2CEfQv9qmOtBa8SDjTANX2blbJw/ktJjpr9rLh+XNRu67QU8GbSqgwutS8bVF1Kp4UgyO9ihzS
xRjpoyL4NLYNlcoXVRHqC596Z+SQ7kdCX0SNwVi2LoyZhL80xjfStu3KKzocEg7i85FsTqSwZhiZ
xOKhse2/FyVnnsErgooaep0jUurToNiDPJpDzrMLI6IcNtEU11nxaX25QZlx2t7oQLXnaqi94EM4
kAuqQPo2EoBUWh9viuCYsmjhz5ueA5r8j++5/xQJGk22x0GEdpeOQdrxIwH2/2k1hMozVY2mSy76
WX7W6UY/vui/dDssZsyZiHnZ8bpaD2WpJG2elYe8bIe4aGJSh99kEIpsjsZ+L+X13PDYBPus1WR1
UVwh6vshp8CDkG3A13HGOVdTYchMqbdoETGJK2eUh6rTXAtheDPdPickXjNtRp7b92h4uavFWJ8f
M2VfY4ETH92LdS/2+5gDABk0E9Ljg9XD3gGGDE1pSaKD6bCPVAh08AP1YIEsJ9sTJ2//cOTh/Mlv
S0BmO9qSUbebYOOGlLmooYOjpRPQhLO9FwPLz8zs+A25L55ox1lbSJlPMkxj5Sd7D5+Gb25tCEwB
gHzmH70iYgQDmS56FA5Yg7ManNXyx4DPFJU+Vh4X44xvZz3/dKoQIDfl61p3vMzA4nPt6fRg4GyC
VXwNotrHT8IzTSG6Jb26f3e/Q5C2fPkgBjYxErA4qm2zUNWdDeWOBdWcOtOll5fjEAo28itibwUs
teg4sOqxOeojFGpnSjLp1Dj7ap9opT8gz9+XKcKcoz5kmW3RpMFAfA/Y4uP8OCLrk+gt4w1EY4c+
fhA+EdJagqh9YBFm10ga+hcSPmdigyGeUzCQ5AhDg5JunijUlLxJhGbOSetBfk/VBFAmsSCgDbv2
ID+hRGxbpR6wJSSv7LV+mgJh2voMLcbe2O5vM5eWj9ZMtXV/B8MZC84dqdlqX7q7BFSMcT/YTrST
vyDzSbVYHXRchMPo6fyEURDRINCKt71nr0Fx3ARW01XKL7AAPTC8qUhH9I5MoWWkpmidiCQecXrM
MuDR7KJSYJrZ7+7kLMP4+2baV8Bm+wGR2SriTQmpz/GeLpGiuJKivIdysywAp3oFsYs7t2XVIg/9
RtteLCGQmL89UNBrw0xcEY3dXu/YV4YNdvxsLj6WFU2+zhX+Z0emZrta1oBEeDO5Hl5bQWpkeqaA
dBuZmUmjV9r/2ubhx1hapZv8ssDbj1unrsD4o6QFTkqK9IV+5gsTB/W+3WgamDUzNOaPIJ0nuckD
5tmzgDpMnblXL+JxW691tWs6+34gVt2PzMLF4ITJHmmd9PSsMLPV1vimfNsNT4mI9ZoDIrQHmU9I
ZTLkhdRrjMTZzrLQKyFtvf68/pKoJE+2p8ELwZ/g8YA+Tb8yfHyVOsV1eaak3pcY4hkjqpF1axh9
Ie0lc7GuJU1N/Zm2sXTPtXBzzCG0tFpfhaU4e1eDHloEYYQxhele0L2vM9d10RNSXGCHdtT9uW/N
BQQduYuN0O4E1AsuLUphdr3TJeduMb59NkPrG4iquPwHwOydK0cvuAA9qpxeG97ZVv0DFGf7FsyE
HRoGLVXt3Q4iJ+34zN0/KmVhVCYDbHs8hXSFBnNh6Tq+oFNQ1eKWdpx9N7wUeKImummVgRYP9fZ1
nTyzno+sig9nNlk35P8N9Erihj+8PnKECedMYdlthxzQvcoClhWwwlSnwsBVa8x5WWooG6eue63s
CSudRkdPxgz28O4tUzjHOD+SnqaTc7mEQOZnMTjLbSd5I7MYouIJ+BgnOBCEjxXV6qv2/vlC7fLU
cWx3HBg5f/0k7zU/id1gpdKo195MYC3C8JfY0YuiALw8qld3aZ2VSbo1mBrquf0OeZYzH1DZoeYG
PHoLWCxqraBCBeSjuLyBkO7QnRzs7nmrDRsU17Ww+CpOqO79eO08fN+3hxXZOAumOujfeP/ROtdx
bfBQL/pash2R+6xhTSp2HnJ5fSYGGzWi57s7bk18ogS71pRelrmKH/oalHVTRyw1zbNS8Hb4iM5y
pfpuzbvIJZ+F10Oddv/I/VBk1NiaqDikBWazZ2QBrlvLvwwiTUqfIu0GIccD4SVN5EMn+SKCFluU
lSYRkornYRbxicUp+SbYKT+zTpJmdl3jJOZkMS/WDFGgX9TEQXCnBjgS0+E0RuRYDZO4cTlCl/++
rk3tiLeeu3bYNp9gq03QkDzA7OTu55R3aMEbsCcILt32d8y3tCkPEghFdGosGTLtJQehiyZjwWjC
6BcluZkwAitir/2UiEUNz6f5DhrkyPjQYe80QavnStYCJtcVRri6TLHxdDdu7nA9ZlCWELhU1Cj+
v0Edxb9L8i5fRg9NUIelzZRiXLpDFuh1wqepjhHzrP3uHWvhdtckO0IgYgzpOP8qBuhxIdluajjv
mFj1AhQQ4JqXVny3KvkZzAAAI832qIguCAzXjVMyh7JZBSxNi6HjKGMaqwTa6lXAcUOm6+gZTg3g
cYxllZK13qu/ZPfGT3Npst8D0FptRRyiV99P75O8ISFBJTKQUag93wVQM6WHlZ4UsIN5bf6YREq7
pyCRc0OwYhRW9MpcnJZ1NsStZejfJ92LHLTLgA0z6sgssbBr1iNmYmxZKfcxWyO0BVuntghJwCfQ
ajP7ACs4eWYCmvBXxp/bUj+n4Ake7TpRXpa0GdgHLdYv1uV7O3odYY8pq3Ns3kovje487l9QIOcg
jZkFnVGqesPBX01uHOYLuRGV/yzyDCCllYR6BhDHsXysp9pW+ABKdgXkOk824XGikU3BpzpC2BOv
of5JnGnqt8UysfuaAWAA01w4izZtX9NpDpFfUXFUl/FDN3RrfqZAHapeDXPm3U2B8TJc6wS0nbfh
t1ywq4/BShC+jNosulb+Ol2JPV3gnM42E2Ghj8yzdsqxjuKoCiPeUQeWVLNylizi/rGxUq61w2Dr
c1VAOH3+5ZVQS2y67bEEJmAm/WGSUQoX/xvsbODypDNjSriQDTBz25uKI0otDA2iGgPBYktVS2Xi
EygdtlNcbd04teM1Ak9zM9BmWnozLiBUP3Td2bD2I8f21UI0+CsBUoj+jTofnoRUSwYWpii1frH2
bCgFYXNavi9Wym1oJXBJM6iangm8jbIAjvVZlKjRgQ8xFUVVD/uyBtCW19MmRRxjgGIEkploupT/
I8HQbjaLiq727VHBjx+nx7Z+g5ATy3DrTl6Hrp74lsiyGK5U/X0EgJ3FKdFFyEnbSCmvnZwXlVGs
wgnmwRW0bvuJebvgEWztcXpOdIv9boEMXDsxrIWG4nGMH4FNME7Z8/akShonJWhRMIfiFYYd2sb/
zF/YEZ+wmA7KgG0DuaEWtU1PtctO7S+gpnm1cwrSwNbBugLxgmS+yMcJ7tAWW10c81tDNJLRBeDT
/TfNTy9kWOV3N0XAYjxWmZqO3lOkdFeOFnIykgJLCUCe68bSy7xmYJ1WxTpGvIWq3KlAuPuC2bDI
YdLNWIE6qXdmy+ZLBQnEZC5UIEBI5o41vrVHIwacwLJbZIL3E6O1r2gKxV4mFFVZRGjNqtDBLYQi
bDqs8iAnv/VEIyvv1TjCKNY+NmijFFvOyyWwM+aYoQRY/5zm9XofacFH8hpLlNIWAqxH1WFCG23e
oMPf+S7DsifP/MJyyyNav489tg/i7FP8o3d/6WT8asBApJgYp+rAnuYrHSKUHBYA1IGGdboNv2Ps
i8pVGEcxwVumqwUszImfv6ii/3i42rA5C4jEnf6RafmcHdDEeTWltmUEdhDvD+w6Yk5+i2ZwY3FG
gOeqMWr2JT6vZc0QtyunULiEvudhf5U2jzCNnxzuWRYW/zH0Xibky037ka969l/lcs19N3WWM7r/
qKj8uZQWmKmZWKKIkA7nYghzoviEhIxTtuvUUF9/2ydCbCDAyKF6SeBvpH0vHjLOjl/MvIV6emO7
XaVU2wblK4x9dAGyMqRAAJt2teEJ7UEqKcXuUDGz1z3jrX20YPKsMJ636s73aSj6zlO6OfV7hUIB
MyT+b/HGQ6k5LX6v+ESbdDcRS4mxJPghPPF3nne4zD9Ekj1M1Q3hi4WD6SFPeOk+QeO9EuomQxOb
pKwUGvO8gFKNbntDUr90ur/6Q/NA2FygT+QJ2oFQmTlk/xzp/Drt/mC1FDX8M1WcQBKXBvHvrmBi
L/8crnqj88jLrXwpoMMdb8Jui/H+yFD7TR2Suv8LJmPpCgw7nVqiC9w/6Gz2n7WwwsMqpi47U2AT
JyyoPqJM1JiMSNLebY3zdvUEJL2aDGRGUvqczd0Jsc2sMR1aPPd/v1CSrHnblwCZEWLpHbkuLt1W
4X6g9ePe7iX/AAbvm5jeLjXUEIE2G+Ni8euvZ3/TqyN7DnbTyKYvM/05gPCAm+mcQiMY5DjyADQA
Zl0ukhD9DusWFeh9GC/Rw6cz2dUY5J40fhTvxD42eNX3FRi+8b+yIFkTjBsqwObY7tGJiMN1lAa6
aY0+7DjLzn6yY8BxD2u9fKXTERunt8xSSYHVU7Iexi26VtbKiQ/auDArHeTli2cubebKT6Mso4Kk
GWv99vRVcjU8s9iIysV35j5BdBaVIk6J5Vu5NVpn680/asCQ+WUPUfRNc5xVCD/8QJxE1gqJmCZG
sudpVRPsZRCKVxSWd3PMerfsMcKQw7YZR9BMGKc90S2smwZ8DI0CXxwRZh0/3wGEFXgTO96yQE6X
YdUEgLeCgdZLEdD1nwsaJwoP4yk99EuUqvobwtOM8/FEhMdMn9VvMaCXlQnCr5GqcNRHXdWYgR1p
fu5QJUhKkmGBPVRYEHKTmu6aK79AQxwPxE2VbPoqyamGKKFk8XkibqNxJj4d4PuedzNc7f/M9hL9
SDZtDTmHKFLMXmStj+XJrJNncSRkoIPzZmboTWawUIpkV3+DH981eth2sFQh6GMV/exqhhgqnsDM
k0rlFFZCH6DFFXwX7EBqGcc9yFde9LwWqP+h6kAb4G1VZ1piZSEB+5u/6s5yOHqxZqHkkTJpCSPK
Ce2Y95B0FFejUEmcD2oYusMT3fuA0PvICOeLAadW0Np/+poAGdg8MRfapM6unB0feldZlsPal2zo
dunfd3hgq3HJk826JYJ9u8W5UwtdthgDVZnF8T5d0WmCMo+nf0xcDsG/iCRM5cWuw0mx/kgMaa0w
WR0eQHJxevhz3MntxkPLHonsIW97brxWPP2Ym0Fr3sNbGLGygrbVL6VASnYpKfkCSaBHh9KQjTc5
IDQQOZr2tB6QRd1nXNv+v7aGFDoLRCChZJ9BctSqd75/QbJT6qcKge6qWpHQyZMhqy2OKgDvyULB
THQGNyAU+X5Zu6ShYDjVgvhrgu13AOd2OJ2XyK6bE49ON6RqSBEg4kgOQghJE+x1hFlEfTM5qXag
y/dT22qYHfqYaApT3yvfhundyuVX6gXrIhDuxMAOI2bRns+3DHtvATzjfamG7+GuGwzzbYYK0dd0
XyiTQ6CZNbQFEoGP19aM4+tNRxHwptyRsn6gW4yvDC4SRDO3Wu1ok2et/6hXe9buatsHxktBbC17
7nI4XYNLlYBs1DMDN1nEzkz5SPku347QGwhc7TveefZSaT80jDU7ZQJLbhy4WHF39hJ0TakQ6D3b
EA9NHZf9BIJ0O6CaoYueRWZBi2fthE/UHoglvdO4AypfRnZwOS2haKi7V4knEidgr+UeWIwjaWyO
xSi0TCAdnzik+Xp6EAkMruiirJWKcZ3PTbh4oWjqMaPiXEMrIhesfTDxCfsyuxEucvO24ZopHKbw
9f1DjyOwJd9Zop7S32MQ3ajELGv6G19IGItY0ZwQDAyJ3aGPPsk+Budpb94r7RKIW4U21gAqjHRt
s7THhS9sU7Rm1YEyl3f151NR6zQePHR0OWfcYPLObeYVm8FFlH3U0dm8I89/vJUcARe5LK+2p/fB
dA5tIfyIhABCp1WUu7WJAN9+MBazSK1MnJV1aGb3ZEaJd3u00uamvoBdIhkLpT5Nrf7eqdvZtZYf
OkP6MgX2upK5jaBjCCpPBF6BL3eIpnb8BcOvp7necWaMaQVe4hn8dZtQYNUOPVulI2/hnyhJRMQQ
ge6V4qxl2kRWPJlEM8V/o3kdnk1dxEs/36m2HyScYwWvFOCLY7RaS/ydTbCrMqqhymMAk9U+Gr/L
oj1CvATMVVcMphiTLTzJaq8v9XhiDY1TH2jPtJ6N279x8q4glaVW8vv3uXc1J36XUObhUEKH/qsZ
A8l2u1Bai7Yher4hBsWw0GJLPW/iiXkWgut2nZc3czVGv6H+lOyTEYq30YPBu/6Cmkl0Ih8QhS2N
OZYDQu/73IK5Z/zsPnD72zML0tnouHehWH2GS1h9Eh+0ZYF0SFSfL9pQzZAok0jxChiU+W+WsPLk
b/hla3lj1WztvsB59ETA94TUNOGnFFNex8xnhErA14Jn1ln4hYYdNmp0i1VC2KehBDP/BWVFh7ho
MDfvMKLdsFliRUOJRM+ySYGTaiAhaTyJvFyZDXiqVJ9LAUUDVVKx/PY70Ke7wbxwUc9VLtnMoL/e
ZCSOthBHszjp2itoQCcJXlD/1erIw6Eol02EdR3fYmfEakaJPRevOs9jQJ5ynIUdGE1hyoC056dM
Gr3ir1EKN2Sq2e431/CL7Y2S2U3T/WAKfppRrrcSv6o7nV+v7/D+newDoszKYI5MSmZnwFGtcjW+
vCrXt90dHnQWi7rtpXASN8z/JROPAiDLfXqCb8hzqHEBxZ/ta7ywt3VKQACiV9pwSaoHqF4AKds2
1QlUy1H6f+SOhLy+k5hxmuyfduqDbe0jUsaCWtKBSWtzRUZV6CH7FhArdylhqMLFbzMKyBqIHNUD
ubJvSDRrHmEd+bbDFzBmmxJUhPiGlsZfVlPZvP+NHj4LWXQFGMDRQcn3BUJJHZQEeO6q7LGiKOGC
R89qXq1XRFEnXJVSHTxgM1+5KXCicR66iVA19kRRpgjpp7jiliqs5qd9oQK9qz51WLKQ5p/11GJO
7MtpuEwahS+lMNYS/L0jjFfbltdBpvfClkOJtCV6g8oW6l9+QlF++VF9+n8GGN0ggQ1RAUAau+RT
Q5Uvi2Z6LOK84eQK+W7CFE0Op8hiuhnbh+Fzs/6PRFeZKG+orQhrwaoIVMHjrKvYzzfE56OYbYDr
k3K7ZsXZXuTINubtdv6nwpHZH9PWDb+RJmBGgPUsFw3G23BXBnegDfnyEchfGMdFH+yEsXuf+2SV
Hkq8yavGyAqBnWjJ8ho15Hx17UmKXZCWg6kkpze3NZ5qXRS9ch2h+3v16Aw3NUt0uR5ardqzoscg
pi4ryv+IRsTAcD3rbsGOfOsf1neHOFUjBCHhb0Zgi+63k5aXo35ip4TgIbWztvOtM2Iq+t85hr1h
GCKMFzwmKry8eMFVOTFBbpvVwa/TnxEz5nW3PVtWxK88nVCFpT4Td59gWRR3Gxb2+KFv2P6JC2aX
RzjP2dxoJhd+KhfPz9KXgsgAgCvvu1WDlVZ89cW31+xLBkzgnrsbIPxAqxGWVm//FZJYAhsQrwUC
tv4Na7LycXOxHB4Q0jvsu1H7h0vtkhswPpIwuAOBiAaWoC0Es5LxvXHuS3uMhov+f+blcA01oyEu
/nAi4Nbpv+xKC1mjGJGliy+tA20TiFlxw3uJqYn3ZRj8yMcKCCaoyG+FG7xsXuARH7URX40O1b0u
Xhe+PLBdVb7eO4Gi/XYrgKJRDxRXPx9gj4Qct1GBOrRzitiSxaLBC3gvSGpnoj/zdA7DB9raIc9i
EjZ8y9sY6M8TpIV+dh0CbBcuL+IvEaptcxgUJ/lcDmxe/knbshwec5eiQeYJ1czZ7+LjAJWphL++
c+qLeUB1Ne+ZZ3dj4KxHtCGtX5a8Tx6WAakQ7rzQFuu5xpPzlSQVEtscVZcqz4pA/liyZUDEUaT+
ndT37iY4xmS2b9BwL6itcJfjawIufktz1eaD5L1PrfGphY9kzu9N4tvKSxktde6ZvDW1vHN9VWBA
HWqgYOqBRkyCpKn9AHQLiXfhe9uwMhi7kFBGeDg5zewfB4rvWebypLtPxxPDESvU6ciosE408XnN
dhEkcPsGFo/FqZwJJffJqE1YPIyQ5uZTDkE99exXG85FzvyHowQBReoWYPR3ePdpEyuyT8lB0hmL
LgnvgwqaRsmysoRX1qoluhdAt9Oe2Jq4AjvezbJ6L33BVf2ks5NhNm94i4DUfSKbeSEERUkvBIX2
zTdZAt9L3JjREftp7VG+Rc0s2AXNHPgBjo6O4T6ZiY4i5gKSyrj0hW0ixyxZBOiW1wNtmvE/9jFp
ztnR21qPA7/34sth3CJsF/u50PB2ByRX3+dCnBiPMyByzR4AqErLnezCYhvm/q76/wtw1bQqNn3a
0GFCgc5rLsxAbRfHyjqQnRdjkw/1m13BruloK5Rxk1TXmF/dXOroeCd3elkyuXd8SZWSJ0tvo79L
i0Ct81p2C1pCjNFzxd9VW03YosU8qsYN0lwN8TTh71vg+amyVMsGlotbhe57MHr/Bi0xH/24fiOM
ysAD+/fuceZu0gH8ZTTrEGURsi/Nby/DWbWH0bfzDy1Mku2MXRjcgKI2vVI1xHyb2fp1lZ8ccNYV
95rpmCtMzM/HFUm8xd5g9nJFWw2Acagd4q7ElPq7EPhGl0L8F/uyYzGnXRvuFMhv0QSp1Wy8dVjk
vDdujC4zkOZsZCx09Mp3s5b1RJG84z/Llfkf+52tsw5lm4qSQC/uVeSVlJkkSVrsbnSF6er7Nh0o
/2YUIFqj+J3NLYNJkL3hDTpYDL7bxGfqNwhf+0vamS8vsqhh9bmV2DUPYKcdblMGAzrTOcsMX/DU
ezbJxUXoaVTWy+ENDeEIl82jeA7epkIMo832Bgm4s0gbTsnrAlC31mU0pYnK2dTlbtvyqpVNmVqF
Z3r2FBm01ZpqjJbgfMChFv7v87pluYVR9Bv5laeW8mLy/VsKe8ssdVBB4TVkwj2777pU32mHm1Sv
xF68SIk40n7zO9JrxiDwM5Ar6kUrZCLxxmykT5MS+YW4qgzhGp8HfhIihee5THLMbs3EliVPhWU5
G1WNKkF6iw4EAhwjdNMh2/AQeUcCafC8lzIUqIc0u87rxbSSef6wLcGa+V4ZB8J6Ro66C9/T/VVW
1OJB0t3UQWNJz3Nxny6rBNRdVyynhmFWB5oo8T+4Np7WkcmIlNZbR3M9IJkD5CyDzh1izkzJzi4e
AzSn5K/cDwYaW0H+CxFsyJhRC/fC8RcEL7sHZY/kabcSCzL9aOoVtGTtUDxRUyMzeKmDUA6KsTOP
X3tpis0xd9Wd6CmWEP4RdRegERbl6OQ9aFOmSvaIqxKKD13CA+/gux7mCkTx2zq9TUILxdYby+It
WgnZaSjv9SSsKjVjCe3XJKIkLQ2jI0OWZu43VhZifZLkeEuh02nSnevdWyKhtpj6ATJP/7Wp2KCx
zG/mxejuyEg+gFifNj6ldDOSj33hW7C1GYN94QYWn/vv+G9VcOvTp0TA4nZCN8zgJJShSKk5TIk3
vKYMwI+F1TA098GGCN4CyHyt1RR+DSM+tz+HscoOAHfhzsznKUHHnf3vXfkDTBjyHeYgoax/TX0M
ZOe3rbox4agUlaw9N9L7o+6cRnKYfo0/HJFA8uUjj/ASLZXF6tpWHOk1LJZuZXS179+x2gqJPoXi
qWZsS91AFvqOljq87dzar2UqIwqYs/ru3yeaqsB3JYcBJtxvg38Zf/x2Wy1ZVoTeIpIPe3qHxMeY
6jkHzeVZDwSyX8vZDYIUj9pAGRrS29m1MjeD4jV7iNWxIbHYu+bu5VoQ5tRWR1svEq9WyjeMa2cC
CTv13lL9FLY1KD639KMPO53EjnTC0ChHM3jNC54wq6cprUQuZB3eFhmCDpfR4ODcWoBMF1W9MCjN
aoF0JqxuF2U4PSafdPB0Jr3AojNlsoO9CQYTv8PLI2c4ovg3/B3wflXH27toUxh6dkgrx9y24mT2
nRJ30d1S8xlfiUdT6Rb4gF5SP+vkER161ezXEwXX0NU1H/9J3ErarEuZGOeqRFp6HVrfWavXAQNQ
dBA9GhlDUSIlYuYl8ypt4X4yfHxngZFvWMskQndLHBMmRAsaH7poPQvKUJ0lHm3FlcEq9N+Z3aDH
JFfDhdonWbXmVNa9M8R2Njx5VQuU1gb6l5v5McisAxYKFuRL/u/H1prLM3q0bzPQr3DMCRQVwRoN
Mi+i2AwTzJYFFZYM5Prh/4NhvOi7U7xLGuZ1KlSwBLZD13lPbzGQgZ67Dr1a2Eb1hlg3O1171Lsb
zMwS+71i+mDxaPO+qzHO0CPt6JjRMlvcDjlsBRoUeOP82nhG6M36XQyj9yHiotTSgdTPTDDFysrp
X19sniIsWkG/k40uRu15O9cfVkkgKj8bvM4/T77nom+dhATz8axbwPSIHuD/MLWRVlBhPwWtUIGX
ZDbH0TswRtwnX8SC0JroZWfNE6alwbQAk+Ny8eZw7XJ57wdaAfXqoMvhSpX2xbH8P+s6npoFLrO8
wPmQOiHHXGzeO1d2ylsXuwzU9iRFZR0QfoNSi4E0A2nA1HL+RrZOMuflU5tW/VG4MoQIl9cWZJmZ
QTvDQa6EljeA2VcQrioO5f4x3fsOS3V4fStip81CuZdXe1BStbsGuD+9kEngLguZLp2WWujAWeKl
mTyLPzEBQfcRODoIA7nuKQfG4tnGAOyjBKbqXxe9pKxR8vnpUTOuWxCHExhc56HsSTrydQm5mTSK
NysncuxfX6gbY9VMb9LqrYy7/bdGmCCzIkY/w4xOj2YPFgQXZAAisZGvfJbbLQPExxYxnAup49+6
ZcJUyuMGANDcmeAgdoK9dD0U9ozRVu8T/TldCmi2BJfOxsZMGT0odL0FKmVFrEH+wylzciL55PDo
HE6s1B/DjkAj9VZEbP3AkvY/95D2oDTF0nU6eI+mmDkIGCMnSIm3av61CHvvH0EQNgrQ1ruJ3HUS
iJANErKYVnyqb2126tHSPvQRc2I5l4caUQu5buJtN/+smN9P7SqMGz5xbNnZJCeZQNcDQHRc875X
tL3K9SZfIPHmFttM2HDpxbWrkrCkL72eLOlkskEUbCPqZQIuycTrhOGpIZ5QQZJLIKmSAm9/Pv9g
nrniyjerEk0a/gBFFQ0sQOSJToIjoy1H7QyvxIianCq2GjdsCreI0K9t74rvbPkhoWwYMUvlZZCu
ojK4JxlUmjq+47u3e8mP1dj9HFyfId1Vqm+/756EXR65zh2bLw+NMg1ZThxKU1DJQIVxA0GhrutG
WUseZ5/nGMoAafvzkGY/bAkO3ZlPmIMmrmkXvE7tj8MK922hBgogFVogIdN7nRfvwfmJuHHED1Ha
aWWjIrNcGrDgMRZEOyRkTS3dh0kE7ObQw2mDCe5HCMBkWl1zbbZeBuX1oYHnfxSmI506tmmnYaBG
/0bFR/cmYoDG0ctm0Chulmo6wW4EjdUtuetbSbhMAk4bUyu4X+SoJYs5EN7Z1RQGNVhAcnqDbi+5
tc3zOqtfDWobpI4Sm6vBcKCLYrFv0DUsHK/eMVJS+pg+SZmG5I8FTt3XoSAhSRD7oqw+W1k9pVoK
ii0PcqR3l5fkHuUKWYtmWXoQrFXg/YhWPvEPkYwr97H5XCONw9lRA8gkhJDR4s7/IdUemCnp4Rh3
aErI7nP34QLxv9+PwnRtNgVWIFVX6JYrckGgVE7SUqS8kL8B1IUOUGmLtn+u3cX8Rp/l8C7uqHOz
EOOcwgrAh+OIIUiEodqsdecsZQCgyAI5Cv7Fx4rnFqFSgijBmU2Lf56lTFJHnA3DVhUu8kXkZR3J
S72xQBcGWgGhql+wd78ef9NzBXprpDt43wPfvwkDUqMzpgcPmRJbkPgDtJ4LyOXG5XI1wHHGWeUg
N/1Ers9RVaQr9oWzruzFDaEGXcOOj/GK0tgU86ng6Do8PnXxb9C6P11bgxpdFxzPFmIYJwujeaXj
JvuZC7CAdJkEDXmjePE1Q0Tu5KjY1AaPWLu+fHqtSmyHp+uhFnad+LRzOqSdnTbT6VqKJW652kt4
RDEPrBqJjmDM6XHvy8lLndnroSqCmQIY5JNLmrrASc2grap6iuVRpcPBMrdX4nYXz/WqzODKHKVR
UERz3cqIHcwy16rZrgQKds9b4u624nzog0DbGFaDF0pKfsXS0NjkR0nRrgKpICucTMUntbGX0DzJ
Ev4981PtuEwuT2yrzySs+myari5e3h2voPU1drrq8MpI2DY9pTHlu8F+pxq43pzmRUved/P/qh8K
YpnWdCUNaH7iaCc/FEFmATOmHmiYxPYlUAx5MXhrFpLBDAdgpu9muyjhSWqkv41P1ichpmQ/LgJz
jxA/KyML3e4zQbMJ6xnAAvQfqzk2UEjXW5qccA/H8z8DhpZ2NfpSAsTWSt9lwzH2+3XmvG3dhZCC
2e5YcPJ+MHITXeis9ut6/gDXAxTI+QLErMtI9Tw/pefXB8XNKpTgNfV3+5w2wHsy7bGzEOc0jQf4
Di/3D14Xq1Y2T9gBDC/KDgJYiJSu6UreGnjh7j2JfZAH7GT1WMzMVSBYvQOx81chsxq+W1jeGV9l
cT0KFJs1S5r7Quk2tcrCEbzd9TdB5HlPtHFolqN2E0voKBaigLu4SNWqyJ4O6tZs/HgSSIGtQsij
LYXtJaGV2ZBGw1fhnHyE97vOzShI8NjOXSW9aL5/HoE87GB/bc9gnMAfSt95NoMWNnm1WSvvIsgI
DoSyTmFuEU8+Jt2U++ZUSfOGCT1QclMJaxtd3Wntu88D235tP3ijclsBkBFLtUMMIiaWkBbE+EQW
zLLSoea6u6ZbQx/nfzppq4q43VuKNh9V/DrguN0nXeRmlJc27AxR0U1+mGMELjFTuZRilQtSNY73
eSidYp9f2PQ3TzN5/MbbjX3h0QkZsGO8J7MWlJJOZQkOuxvGvqGuah9C+gOCZq0I+xF8xk933DWn
DbwRYkD/Q6lSdkyTQ1MmONIMfsc6edz/pUwHsQnDJ2cj11qJdJmL/0LabCZIHs5CjCC+75S5p6Ll
U0Bp8GLKG/vqzVQa7eilIGCuCS2dRUPPzYg6ewSZqaZ5iW74j6/Uhx+F6qGDg55ddyq6f7Fnrqf6
1pL1z4ZjkXlIhy9ngDu/vbZmxRlxcCWANmy2Jh+gMgp8HHYK/V69abR+b2t5BOoT6gUP0GkozwHp
RuWjsMskWAjeX57j+nmjN8vz+J1MaiNniLKjU/hGvJIGDZnLaPmt+Wo29HmwGPfykE/nfpMaZrpr
D4FssHj4/367QXgziIR12oD1WtgCi7+o7m8yhmqbxEDxVMTEEZehZmZGjxwg2hWHiPxG3B4H+atg
v2odY5dKHXPkZVZGD4D/CgcaDaRCINZXMahmCRj2nKJCrscs5bhLxif7CIxF8a+JUy4CQZC1DU3Q
FWXAoDpLjphFZJ7f4kZrkAqyKtKFAkSDME8C34QgQ+e2FxtZAR3LMU6KYRjURLBGPJMJ+m68ShtX
L+BoEuaXVZwr6q7D5mUbO9vDgNygRJfmaJ/TlVJNnZ1rmC7a1JDYyMVYSBgV8rdi/WcyMOKlHTVB
+1iQnPUe3lRr8aaE1mSyt+ZFxN2hb8dOO3gcyQYv4C5N74AcKyl8RsOzF0zb4imvwzNkC4pWf1M2
VbfUhdkiCR0tMNc0PElzcjUm7VbqnkK6GbQ5TLuTuDZqQxTz7sBKpy677LGTFaglb+0u5oj9D8av
ym4hW0lp1THW6R9exshFWbM/0JHm2hrikw46acPBJxvM2cUFlcrWd8xIm6V2wt61IoiI/YKbBHop
6Q6AQxqe3SzjX85/B1VLUX60zNXzz2XYoBf47BaLKlG2lMEw8nZZkWmm4HMxGWjk+XNRT5Feavnj
bCDqnD9/HLeOa5kSBE4gk6MnMYTAL6yQIpiKG94VRWCC9h75bE1jEzDjsBwF0+JQox8EaA7yULsP
KmVMN0JshiXSzZqJgZtcWa9uVUCQHd3jZADzwY4BxEjYOluluhSWHWt9uKozrv8edrUDB/zAHk1m
kOlgxxhruVZjgdc0goVesWRuVwXhwiXKENF0Bc79w5NcworEVEOrv2WF8P3HCivpjgnMj/xrO3Gw
cYXjh4+VuL+/U2s2HjqCjh+9a+zhuSPjPqRTkybwk1xSgoDuXbXdtyAcwIYyhvi7EeR0LWHRrThl
Syysp43arp3gjpOb8Y9zIkOe5PJozgXzXRTl/P+t8fyFCrcVC0aMMlMNua0rDae+XfUkQ9rNKBYn
tctU1FOGsApu79cxI/iuatMvZvWtRgIA6AmzKUcDkREiV0rKaSOgU2+Jp8+GMcOvq+o8UXXiXxxt
D1rnwGqg8aUDfy/RIoSWe6ob48y/kkrjmcSYxkob3XyRFbcmIJ9I0AXf7eFRcy68p1X1urNP4VTb
Z7oEleUrIlS3dLccc4DqCFmUCKDeSlYows5DEIjASn/DqgdRHIYEHxTv+Mcp1v1eZTC0f3lhBIfH
l1r1Y541uUHOHTniEZrX22rfwBZKcMcyAhk+woR0t1RjQAoq6vKAY9VdhmzakUWjzCd0P0Pb46Wh
yJfUMNpG2XjfR3La/sQoCpf2SZFQ9fCzHfWFUCqrXHU2HmAfbbaUOkMeqXVnjrSstxTLhPzAZWZH
FsCyO4gr6UMfS1/UnCc8yiT4VGsUUW9wCJ1LBUa2i8HzoqwQvSyNG02BPdp2J35xTkcWpEOD2xa6
TJrU2kjLdPn0Lz2NKnegrw+eGF96kTGVNluFoxX8L+7XkGlorWDhtynAWR/ViGdl/6hVBWCKm6+0
RjOz2DMb/rF6EA68RlmoAsLgRXRtbsMqmD7oAaTakwRjpiRGTx1KVjj4lqIT5VexvW9qmLRLFQP+
9boMjB/rHea7Rhgt3L5okmhrNinf7s5JaDMlxdQW3K637R468DvxsWPoWJQ6kVoang6uX6Ol/G0h
s3CQN6sn7v3GnrOfdsycGUykOa21KNMnW9XhK7X7Iu8fqk4SPg3MWtbxIuJpowIcUKs46XAaC8UU
80Wkeia0jyPKKlHt/jthYiNBbMfeOHgTXYlRGgFJWwHpIEqnM5BHM4v3WnDH1qbAyhph2lW4J9nZ
2FGWrKzsHM0R9A9qUtigCkR8hejCdiCGc00teUS8RpuA0zRGffnTUza6kJ4JFr+QuAHB2TU1K7DN
DjVDVG8+WinUKIPFf0ksmi4Ota7z2ictdHgR0ORXM4FGnydPhvw0lwFhg5VWa5WVBmrQTmZZ5wdO
qJc/4s+DL9cfwvVimucnCuasXSrCmcd9z8YWdRiwr6UB6mfLwXDlc77Y7GEOBr6AqgKWfVG1HeOz
yHYSnqagDvzQN2gwdmpUB1JX/ZkCRjWzFOwu5+LR6dqMtQ17dXiuHoCRE8TtSdgf2KILAh9O/wOi
JlUzawitRjbCW1ESvMbATNOulDCaNlUSXUW5uT/3JT4PS33d18rWq9ls4Pj6RkMOjqQcwEORaBIu
mx63GgrQBkuJF+TRr+bjj/6rszD8JW6U4vFQhDteepVf11K9Ha1CiDdwsik+HHS9c7mSXj2Z7CNG
aMgXTxjXUK2FIHourp9wn/Xkkmvs2/vWctS9jNu7cuCFATT8RsPxqL7vXD2rXLN8yr9/Ze6LwSEp
xp1uuyIl/faLSdq2goRgspi6w29dqYnU3cH42grqlhymh5EbzLRBKmat2QXm3Jp4kKcCXhImQdHW
bNuYXRDZ+WsFXGpYgdg0OjIIa231jfcekEWnXhBQmcmBIERIlLRJv5YeZjQbON9F4DNcZNSNsFOo
g1XZQTgXc+XfSnQIvqo9bk7HD/8CqnTfChJENhxmJHfgxJVu8fheuOZd1XlCugz1KbR6JSo+Ltwn
v8bUrQ7YwiSFeDZ+5kdQN27zcqYwwsoB7Bt5KJ4Z1jBLUDz7BxgfQ3DISePOPNUaUiBCh0VSyvR1
7U1C5yTr4/Lt+8C7p1hXBCCqy8CCtCIPw0Vg8rzmotiGL3T+rskPRuWhOgbTeoB+LiCbDRySwA2H
5SeDDYLIxwzH6XJHfxa0N2B+PWGNLQ5nx+/FoJ/b7R7fdsiED+/FX40nAJvz92vgaCX5T/e4K5AT
yjuh3BiVeX2WHG9nVT8G7ImIk1DwlhkaPeNeuhBbeI3s/QELMbNBJDx087OMTd+Fq65krzxFDBo9
Q5vAN0gVlHmaC3bznVGSAzMIiP+4CxCgJiWM93DXvC1G4OiizyqiTpq0BvoJDS+n0ilj6viSPS0b
5wNSg4Ik2qEp8zfMU0ZMb0pQaXRsavOBnaYR26/Gb5h52Zyi41+pdkA+r0CElRJT2NqVOAYCHRNo
npmSG8Nkslpws+7rvveyBkNbGHaAKoMyNRfYG9aJ1go5U2rm7Ze5iDl3EumB10YEPHNNBZKdCrVe
76YQgW7Zh897aR9ky2/xHh9pWsvDKvQSsi9LiTIv/9vECL44G0QGKD2VC/oVvL4sNaVKgk6P8U/R
FIVZZNBY1iFUyfFplvNQDROtjVtVLPiDxZOUf4dHo+UbdZ7ryUoqCU+Efz+3Xss50u3X2gg0RM3d
AvAtdWkhEg6oZDWYy5W53rKFUfCqsE/Gq/Gk4uprK6wlTFvsdpVsBAiqkYPWajhagKjT3HzS7LFM
DKMUq0b0DSqEIja00Cj+GnBBwngoW6ps8NEkFpQfd6cVtIvu2VYCMvYhJvNv6eBXyARMVHMqsydk
jvY8IGkRY0vMN7XLn4hWWCZZjfBQbL6J8u894XAdaM0ThUyYoBDDJj91cyVMn68hA7gAOxKGhBj/
4F0OLgFMZo2BTcSOA3Sjme/9749ESuGojGRNp4KZXwxkcSwt+kej1iLEuyWlhqZzGHHS4FytEYXg
73x2M6IfepGVkJGhwSoe2KLboeebi5cb96ufQqsmZQHYVGLD/REB+gOXUiI4g7LmvAvWNsPLpJA0
dgT5ZbXVZ8UJUvyjUMWdN3i8+9eVydE3U1W233S33rcy0sae7t/aCOJyfHG/q5o3xq1Vt1/er+ua
febZnE4M76R32+jExxdI0RZhOhfTiTY4bYCIHvJP42A/1KmnE76ifVck3IiRax5J9Tw0clk+5u/n
f18kQsT9xV2YIe2LGLuBsrIpXCIj0wnGV5Advv0zgksr9OpI96v14Qm6hGYnNPtHj/yq96HGsIk/
6coRxxyxAx87ZiU52bj00VKyoVAqpkWSOXGVrnAjPMTs2HpofOVoLALioW1ihizW5TUk0kK3BzPv
85A5i+VX5vVKxNOX+bH6O+/hEDdrXA4ISvtlzFgk6+U46nmdSoN6MgfNEiE0Sjwcj1Acm3IdAGlq
3lyaNJVztB1FdyJ45fVB66MpeQhQDcrW7l1ncCeAjivKSi/9ANn8G3EhP+gVE1hFMeuXWqP0JNsj
gb69mXKY9JaCgdIiEr9BsOwqardjkQUOulj1EQ7qmweT/eAmX9YaRC+0JEo4hpMsAgLKf1aMvzlz
96GDZhIUBkKxQes2iKWAfzcJyt1wFqPliuGBTJKtWc07MQmVec+upR+BaHv+PMFDMrlysyROe4hM
PXY5DkPQ3YdNYZVs6Yqdw+QRrg/vQ5OlYxq7Gp8eBrr7ZvGTbN7pF82DJs7CQv65qE17aD5ewWM0
mz1GqyT+Q9VJTYxxIyEr6EvtQsyCb/NnDi/trWvO3RYBpapKkOi9RMQp5mVijxgIu4nq2XllY4I8
ockfOIK7UNIXHFSrhJqgWwLFdxmrbWrBTEE2HG5GpUen1FBaD+0YpUUyQXdmcCL+evPAzGdRcUj3
sBBAm8EvfThov7ynNWm9AGtUY8ZWeasAxJ7V4LixT/3aVwIU+LssgmiJdC23eFo9C2eH0CC0zMTa
D4G2NRKHytIrkpEi1a05I7gqnSDA2D8azOOy23FSBllaEaMV4lpGMHC9jscqJ21C2/CTD8NBSvnI
UxQdIBnpCYC+tE+w18rbAFoNTJRlcGKjvocGVR19VEKyVebgrO6BaOcJP86JHe+yv6OcNAJz47sq
03BkK3yYURS9ojwBNxDGKd1uG41/1LdlCkX9YvmS9oHqn4Brp63DTNjTWmlPCulK57pK6RbNgjN0
qGZ0rqaudNqFYC+czicJ0TmcxhQLD+DbeLvr2gkTGG2V/fSYpu9X1lV5tEcI75pfOVDwC/xStYBc
QRKB5iD6Vn9ehi7vzIyA7a3X0w2M8sb1hLWXv0tQ82e3D/J0d0xC6wrWohtD777uKJ1nVKpkyqNP
H6gVls7JkJi73vfEj0dmMqvjWyw7YgsxDy3xOY2PSN3YgJjP7QfX7qGcSR8lPYB/o3+wK82SoOKp
1xmjlXRDFEa0cIx89L0wXF8Q+J76x5sWr1darriZ0rDjvwzTwzlfPM9/lK6mrCpUT5t5hs6BRL5t
Zb+CL7ktP+R1QgpjtlKoXp9p86vkbtIuE2TstsmXptgEc5RU0Z+l1qusLfx1qOFiDZx0uEQLmdcA
AwJ90qBFKwzH65yEy2DIBfqUD5zvx6XnbquKXeaHAvvXboQBMEk5prblxHvgbqw8J1fj1Uufn6wK
8gfWduWSnE/SJrQFMHQZeR49AXiMqaSWTJU5tJQT8O6zgQZLn06eUSo5VhMq6Qddv+imFAn53MNf
5Y/6+9vfWSPbAqP73EXUyO2dycBWvdn5srcs5DE9f0ne029k+4NWTYhUl0uloegKG0apvjQoNySq
ekypQBI8K/U5j/42O4Q7cdH2ia22Gxilx/vWCIdHPXIE07y0Sa2gpl0sTp6x9hPTRo3u0G0JvNN2
z+8ThCOoAbw6MjNH5adn8QJb/6cyyMAvgnr1lKbKvoJ5zpyWm2zXfeomdLqOesVD7/YqkF6aZBJI
9Pt6OO7I9xprhpsGHrO7xiOWDJ9LFYcYioz84qlT1IWXlWKdgscRNPLaILiZL7o8sN0myiX9dOh8
luzAAzjyPbaXtBH5tN98tA6sGTyZ3gVL7so6ywmtTQwnEkeLjQRDbwPieZX9YYWt6YuQwtUhX3PX
OqqpgxwucbDCiJOIHv8zLcgqjJwwurkpsuHu9gHE3her28odJgDp9E0Jt4p1mkcQYKMd8bsXmjI1
hoBjDNY6pFYodr/YvriOh36w9Z9Wosw99XFOrskZgmeiWMMEbPv2ogLZlENYFs9QbRZ5dbjTU7fq
2lyZYTeut0IaOJvmTfnCJiGrEBwQiX5b+xC53uV7CFDlgC6DU3Al7RX8GX6nT/kZZUrysEBINbiv
GUCDwgQR9cDlSLTqR7Z+r7822HtX3zZM4T62IDPBlNTr/uKv9NGggnRMo8vOHiK9Gl2yUDP33avu
COdn4Gq2W2YnqJ8P96/U3RkLxG41XYqA7pU0zp7V8mwe+Fm06RlCXXDPISeajjp9KuEDblWQT0Zg
MrwG/3E7VhZeBQXvFsTjvY5TOTSVDDNeMHx/XOA1w8Jz6WT+bcsyZgyEtGvgjBR0WjR4ILh2BaP5
TDGXLhS+hBd6IYlpzJ16Fo+KpaEU+CRWJ0uUDBph5uVGWigNjV9JCq/w/EpbnozRTGfmdhAEkKAn
B53BWGZQDRw9S1QFTpQCQe8wyJF5Kq5xRDYadx833ko2K/WkfBxVN7vVW5rDMAMlEFQVpYSRzOlB
8CnHFlfg50CZz9k+GryMQyip31GQFmerBIG+1VFXC6afAHNkrbzX6bcwtncMM1nQyGYjQqWCTKkf
LE8PV7bDjuPZoHtDCRndOjOj2Z1UvC3ZzYh+BUsDVgBWwxg16UgzO0KpuJ6fGBNiFzOTQ4tLlDtK
ql0pwmL6BkCcS1blxsQZ2IkHOCchY9/13PV8DrmPRwt0HFp+H6OK+9rx5yFrwUD4fDnWS1qh4pgU
y8SxlsS+EVkA7ylugFsYcwM/v2WRA5qjuewAlw2T6r9Tnx8iffdh/D8HwCTDDFD4DxLQRfN1WzmK
xksHIbo9AHSsXIW3uYnWenRbjSCqBbD/2+Uvo1YDL6lVHDov4lxSb20Vq87i91DKsCJP22bskfAy
HMPyNrCKaFN5L22lnGJ67gdOMNkVs4ave8ltAhMdeX9xRbIRJjFLxO5d1tTO7vR1s217kIB1EfP5
l86z7torqwyg1W/Dggs0WXEGQtxAKc9fYmujG191Agv9bdJDrQllkwm+uWgmgw954Ax1lW0r0zVZ
SeXfyPWA+ay5dEeMOYnLbMa+jXtVEia3ilcB9hMmJmNFpGroPuWdHh66rXJaGESz/gANkLDAMjOJ
yiXz+QOeE0pe8jBTf2qVa6yeMTi18SI+6BY36Bgvap9Cb9j77P2JTMgWMViNVDBZGK4AH2z5Llaf
/bgUALG7w3QczRLXGpsP+1/fo5ietJUQStkIIjwMh5wo3nwsnyHTW/Xwwh1TjSz5UaJ6LOEHe+ef
SRtNwHnsdEDBMGEodOC6ascZtTbtTRGdpeH1KvVHs1EeZ2qMC4xIWMPACnNKWkbst4kUM+n4NC1l
seXWW/9qLPB0cGRenYfXEhuXLyr9wGDVzw8RQXPYr6WyExvNrYQM++c6vSniM4mTvKfEW359VTVZ
4X+tHpQJq10K4kiptXfq/bBTStqz/t22fQXSl+NYvMDaT7AXRlVuaEsidwIbLhUOpYDKCYWnpo5w
sT1JRbs1z0Yiwl/D7eEq1QhJlTpEy6BdlGhVPCfCt0JD47NLxeNyBqwHUoRQV7czVQG3x4FRT2yD
FehqV7n07TtjLSEISoPxWs4DPMvKBuMK7wFppFinJ3C5oJRy2+jmnO7baL219irgXS+VkjVkJlMJ
Hvlznp7pRMXziVkicSFEVOOVMS6hH/biBLygxOsTv0/ET/5ZMjshysb+04pd6x9pzerTp1XVa5KE
ut4EdRlV7NoB7Kd7vKbOFEJNCIzsq6YiyNEWtlgFILgMDjxygRtYSiW6q84+65y7JHS2NnkcWjyg
lTiQEwAIda40t/HNW2ImcuBcIAm6y5APasxUhsneG6rQfh8/LYxVj55FMWbaEmod/aWsRJO1ZCc2
VIF13K8JGZ3e0pCkuM6aN5YS39kY+Et8qWGt0vUZZrYbCARO1gdZUFI9orkKNuns4PHUO+d5bf1v
8WXSH2rMdbYux1xATGo8BreosNpeLPhwQ8x0NqM8NcisJ1nGT78piBTJG8Elh6jeyh7zFE4cNaQT
ejI6rowXsEWSCMvjanpjoiJ6hQ3pPD2ITE8SOIZwa5snSVcBu6ezlc+ff2YsFhL1wBMqYHzeJMx1
Xg80j/50tlqDBMdtjw4CR84T03tYQn+Ox19sbr0cggF/sSCdqJ4HShemMJ1w7a/mOEYhidDXDN1A
by6i83lGWh+/7VLUJKJ0vX8bneten3xtexd4UCYXWS2gRIXE+7Nz7qYNvIq8kuESgmAQN6pXkUaX
beLB44yYGLQDRkY0K1piiKJV91t6FZBf3N1ns+G+rt+9zMFgBCP58fPFyhaz+fMydISbZgFDK6uw
4725WKpIJwoID008Zat3RhJaDXq0iavC5Sb3otBC826+fm8I/6yKdDLC1BVqhVlUpsS1oFpV0nM+
nmOYFbzxq65eCXGN/yTM4cCGk42bR9OZVYfI7B+ePcNvtNA/Fc/lNoovUwKo5Q7gCjsNMshU5XFE
xcEJSUqbOnHRMmuJ0mHJwI2b+B659noKn6Ym4EMMWbsDe6DX7NoFc4RGxnnXuzkrgWKkGxIKb44Y
gRM/VNtQI9VmabA1MgKqJzbUoxbUDy3qogEpPuZmRxh80WIIDUbJWkB2ws9FBYaTKCBnfmtCK6nt
VYdf3hqFnb17CQG5RfJdaRMCwkLDdRVGvPQzfag6S7cENwIgHHFaVXzEI9ow8yWFi3xEwrowWCSq
MnOuM8CU2/xp4LG0bUN6BCzqmymCO16V9ntRbijt3KcZK/iGs0NFIVxLw7T/1fbZ1YReY6O78cgt
e2LvPASKeJ4H0xhDPCLhwxkfM43pLmU0wgA3LDcNax3wLgF1LDq9yX4clRLfWkmGpFPWKT6k1Slq
lpDi3x+kf280E1434yxIW+vh3n+9U7E3RPDCoWtMB+oZh7sseYy4pK5tFD+RnoKm3tEO7gQzNnd3
zfMMvLl6jG2wmoiR1vXaB715AWHcUMzce91FMcP1nU+d9aBAGJwzpJ8yFM60eDHBa/JtCOAsUS84
b8xHztnAgRLT7GZO2tgJz62CshTTBMn1q+rfrDwF5H+09NzDgPU5XbbzgJAsJRKi6DLmFJFI79zP
UkXJhgP+X0gSph49i6uaFI0PjFuchUiiIrTF7Ryh1pTsJsdgIqZ2Kxg4Fpq4oPvEBuLEO83WLcLo
GqHZ/BLdoDj+WQZOcp0qQdABGTAqUYQ0vCz8fH9BPUhpBuMMuGYdVcvfUl7sgyOhmOc93XmdCerK
oQLr6hJ9LDWYoW/VPgtVB6QvgEL5ncH3rU/quDv7+3yxJTMvv0aXy+FlKJiXzh6r3kvGEpgapS4F
cwkjQUfJrh+S/1y0ByNc7Kx/Xb3rSoQMMyjqaEVnsL3ycn09QqzyIj3PunjJOQN5kTAx7VnIZ8O/
kB5BoqhANiNSZrKZyZnAKZwYwTwhhb0vAqYuE3DjRBr/vMuof+biWn5K+e7gp3EeEFtu+36amR3W
KOkDqwZY0esROq8QXrsURQkgL18VJGtwxO7HNof4eSC3Ai5TzTV62Hv+YU6HUHiyLQVYvB2Qw84f
mIAekhhDhykN21hHrI5Pu1HArt/5iXKBs9jxuqH6gm9P8XuYj4Q6EsFc683tYgDKd/CxjzFpv1n4
a9sDI0TzEJPMXLIkIZLmFmmhEzOiWV9qNOeStjEbQ/ZYnjEdbMs9BLymWy6SpBTGOqIjnGzH32+K
dEjIk3nMJdb7LNCV6Yd4UNfWMFrk7dWJ5euHrhLIQ5aKP4eY1Q+vDiKc+9cYIsP3EZcUfMoBi28P
OFENQZAY9pXeNDP6R6bzAK51Za1daj4tkiA8QdUrE3m0d1KtEiRgFjmiEQ5O3DdJ2L6BP1Y1Vxyn
qn5/eDA76ROA+MiRoRw6x+txta8LFqem60McZrU87xATWM2wvoEW/9Jxhllics6GPMyd3bqRwxqP
k3GTC3ZfBHB5J1hjRVAkMX64w3HGiODVl3LyoSXxFftomtSwqMzx9TKO/+ID+9hTiNqeAHMq4fi4
pWQ6XgAmqRMVcy+RVGqoKMj7K3uF+A2plv3nPwqqNKaw5C7vjus3hhf+61SWRqTeJ0mjCjWygkOn
5IMeioHx+DMWUZct58qEj487zeBhq9T/01768sGmQ5pqMwtpFg/8h6m9FL1pPa0RUKhQDtbTTTxD
5QXwrq3jGGhnZ0lZhe/2fQoabERFUQm89UwddGv+78avBFgr3s3/QgaBTNa8XVaSdnneUTKsq510
V4ifMMzVKFWVIgx9PKSYrJTbKXN0bHphy/5T27oUps1e1+FoHXZ21MPuchw70R2YO1Al+R3sSi2Q
S5hVN26XFfmJ5mrAOexOo/ld1EgaACsaFkgMjjw5nhIyTgkieg2oNVtM7PEWwx8KIOpHsK2rOrR1
HE7IUB+ueAU9Vbeokp2U0rGDyQhKUFJxpKVsLkiXcAYqZ97iBC0B6m7wdB2RYPGx//0I7Fcm/Qd7
CcF5PbsU+LrBA2krXjOYoCIwPqm3BdF+iQ6jOjQb9Vse1YegWkvLzNJvJw7arjPAj6B6JBqhPR/+
WtOH2HEOjD6DfyCPVBgYF1NUduasKszwDdXRrrSg7q+CRKTAnd1SVbQsCGWhfLWTbXoaLVutXUvh
+pV2SMB2CPd/Unbz9Clz0SMwlRhvd/28L43Z0WQ3xHrEaZRAZujMrnXLTtjZW1FsFn3pSVG0pIOp
NrkZS8ui5ZfMd+q9km/0D5royiZnC4wLYnY+bKEGWccn+Ge56VKXuLV6CuCsgJNB6dVml0zbzIGY
fRWTx++SKIp/6/U6OAQpg7a6z4uzmn2n2ENBjzIbx+PUHY62ngIJToYtPa0IK3zJrMkk58aj+xtm
n1nMzaH7d7vl/x9tB2dHYu7J6SmSns9dsn35Yt+/HAf1so5L4PQy010kPE5y+kVDgwJPwWLaxcNh
gZWG/PygHepGzIVjtUnUiTkpLpwRf0JxEQLWcxpC4ifPP7XdV0Gin1wh5jT0emYv6CSFnXRrEDVk
Ir4G6jlWoIODcqKAJf4gGIFD0cr8/ddvqPkIrbgButHdoIcMA6kgXqWeNEk4oclEnbQzcp9Nj4jp
iuXReX29hTSif73CX7+X/Wghfx9rbu2aYMKm42Zw2KZ5RyQzPgdawgS2WdhvG24TnSLGcOHPv4H2
QJjGByzlzh4Mmz34vKbrQ6z1l8GycpKv4MptNVE9cLbKcLPWfnSkFHXYzscm5wq3rwaX0XybiPJD
llzSEb3Lsa00zM+ArZuWfyWunzZkuZUIWLubsPj8XTFQN7zSGt4S3wFc5r+eNfJ0wM6uTF+7jsgO
77QsjnG7Z5DXBFUHOg0mnk9qrejQIg79e/aq1Xg2dbcztAKLR9vWHBX0ErPOCn2eiAzF0scOrAQg
ZPYNdfZHSZTXJLmBXy0jP7GCDgwWXFdrHTubGpqdOJz1LM+nRPl6VPKRR4I8VxxYqbL8AjNkQElU
55bj5qIc/XNxq/9ThgOQgNNpstU8vZEXvFJA0d8VFekCM5WgIEtOP5saZczcSA1ivsdNOgaRPkYO
2atl65TshNe20Ic1aFoX5pnImWp4IaGMYVGigW11i0Dm6IeBVk2LbXg9S/J/Sc/48D+66Kvv7F9a
bKSIAcWQ0dCIm00VLhk9UXwdhCGjx0SmxzXW+3yl/ultW27TGBBvFE6sU5ocxmX4pOIccjRGhZMu
xcox8TRLKfcy3Q0aZC/3rUVyOm1U4PU2m6y3/5sqNCtdmiGSlfUFxuNELMiGv42NN9Byfp37EN1A
gegDA1kixkWTftwbX2AG5c/hfBcCSJPnYRWOlAxj2k7sDhvup6u0TCEHFresAiMu+gzzAi2bSICU
zOVBRC05ggvjAMO5Cec4Aube2XLgTwCm0EUyPRGVhW8f7uzIjAC9a426mgCctNwWSDvgG7c5+0oY
+pOyudCJ6lyKsBFLGv3f6c1SBFW/WailC9g3loXhkpaixDtM4pesv2tpwBx9wC6lilz75yx5fBOS
qAgSOKS/LHHNdKmYV3Rfa+Wfon76tI7XUtme6L/V1CwVox8II9BMQLGKAhd3x3noIAoqiA+5L7sX
Rn4CYCWrDX/LzNBU63v4XmE9Wk0LhOgKsMV/OcOXjYiUe+0cvXlIIN/dcfJv1n1pK5jhEQb7HL2k
WpYcH35Neth8a/A1VdW7sroBq3xaVJwF/qMLm6T0YMA5YM4SF1kX5wM62AGblVHVH7CzqI20JxPU
rhMPQDJACnHRUh8LtyMAxB6X8ywPcOnoDwVBFWpFZdIFhNcOllZ+T56jHW4PzHfM8KDV5x6FkTWD
TeXFmDcJuQgLMcG8MLJrSi5+S1rxugRYHN4JVEtGGMCstkcTSE98gD5Zh62PoWbPafrgjHnrdd1v
v/6RqfyHFOgk1f9PMXjap1yrchUN4DkTXHca8sW9uny+E4cQy4g+3GlOs9hhs437qYMm97xk+PGH
5j8s8QeudK/EnkHDlGh/fNCTibG2FCNieOc33Y6GAWT0WyFbo6NL7Hl2FXKiTlyhM3V2/JLgjRPw
HKgguFI18EE0b4qtgsqe5xd857gFksyqzp1hiPQRT0oTc43e/o6ISe9mSfmyMlGYt+9VekWkgDhn
dwpznBemGed3pWLZ08BNFPRjsePaxfzTwl4plm4BQGj3gWiXDq++gxzibSWFHYHCbEptw5Xpgx/7
qnPGhTAobpnd2ZhpjN2SXGZY9EQtt6LIWQcxdHPe3mhHrbVLHuYBq1eWdsPV+OHr3Fw56nyfco5E
Dw9m1iN8lpOkz3jkQ44tKWVs6ajovfZNqIJF+uS/VOqc5dtv7uuPls5/CVwII26A3lrf+ye/DoHF
uUMxBIVgXCYeFauuoySGuTiAG3Xag4P5z5xtMkpQdsPh0MEN/FeAoxopc5l2fveC0LnHmJy2po4F
Hg9ZUrIqNGO8L6u71PFHW4ZNY/xxZocyVccsqSzDzqGF3zGIMBNHwNjBiEiFPAUoQvKE+ctUrMLy
s6OHZ8gH2GZknHtGY+pnh5u99AwxFwyoe4w4xDEnyBJeZzvgJ1kL7StG9aIQH7V1yNU54ZwjzCVi
gq1fXFwYwNVCPabL6e5JC+uQgcy8FtZg5nhpG5xW/ofdn1bCe1BJWGEDY5s2379mTeN+C/PackaA
jMAuhmMMYS5GObfih+MKNnqgYMvC62t9sBZ/sI5j8AAR3uK+UCfL69CcQFSnTmzgoqE4S5ir0GvH
3uBggirAZzuDzy287iglrH0mxlsv9BagoNm3lYnINwpsGKPDT7bmdPCklHDNcPDA56CrzHq+YcL+
I3tY6NwrbOHb6i67Laayo/6yVmFpt1kJjg6sVPftaQpDwbmKLOLbA7gHB1tCF+OZ0IRmlB1Ve1ZZ
r18gnkOOCi6nj4XaxAhx1ul4ZLnzTSZA4TMXNtApbmS7coUY3FWrrK+Z8BdXGLRavbL/Lln7g9qY
uNcNhchM0LqED8vkscgd1LaTdScLjctSXWhPIUnfVkwfPiSr/oWBhFrGd1zxYKoKY0302Se4GZr7
oivmUs4wm72i1w0aF8t0p0ZU9zHVpa3Ke1wy8t27BT+AZcXsHbVi3F94RKA7cZkHtB3SbIsaxllH
6CiYG+Pl0+9Oo9vQWlFp2DkcAyOk7pH0h4RosVNe7Lxoo8I25gNFtm5ejiFJn5kGWonP+RzXuYZ9
Rop0Lv5YDGJy3AtHTB48cfVdi0xgFoYcoYYgWqAzUyX1WjO9tcU6DP2GOQjMDlQY8/KlJYkr3Uhx
FuZ62CwoTUGkb5inOKc2i7CdHG+oqOWnVr5a2VZoDjBW/ulvSPgXz9/9X4Pvx78Qby+a6XfMKLdS
BkjcCtzqzxqfUMzdusANDla9omaKLHTvjfXITQ562c/LRVzkoPkeRAtQ8WlAyohnD5bTCwfAi83d
Ng6a6K+fK+aMQoi30qIq7QBXU5Hm24M3R0P3IwQ1uXHKzhm1RlF5rQB+jidVosUgL+Sza9XmmPeC
ynqqnpsB6qigFNIyNFag4RMzAlpQBL8GuDhnjOGvPFQ+yp40SRCxhk3odpF6l4/wWZ39KgPDJ7W1
QY+h7uHth1jD+M64fIKvBmccob/Lv+DkzPYsj2Hz/WGVu9YNKpr8nNDCXdwlpr/MAPRakTMK3/ba
FzrPdO3qyAN9q1EqDrmh2Qha7L/HUp9q88H9obqC9S2rj5EMveQtpM1XMAP6qycE4bBAegfmWAmD
40c8cssctgV/46O1fz4frpkICoG7nLK0hKiOpIG2eOIBuRfZ4r846EfFucgAK620JIkGAcPxLZsW
2HY0wqOZpJCgBGnBKpj37m+Lo7K3p1vt+MEwwWAqSe5szSLx8sLedB4yIRhDSaTjh6VqibRW4DHl
U/86cPzeOhClmtn06K26cKe+C1KzJeNa7NI6456FWGukHzvRy6JelIXwlgAL1K7IfRiEweX1CV93
U7IaWmKkik1KcLlnGh0ufaxubZVAwybwNkOXg/YkM9TnJclzxABgoNyiTzmuKDHBT+FIEOTzvP1D
FGF/LnsBhZEjh2OAN65sDxR3DJSkAmBUwId791hjJcVs2flFagW8GDJqqI50V4pRv80ikhUD87tZ
wYRuquHuMnCIz3JTk12iWlBLHkkkFdupOjKy4DUd8VbU4Wl5T8e7zYNRmCEENqngaGkIdEZOTxPF
0f1JiN4ZhNi7KgwPK3K/pGPbhRbofhoSkJfaWXbOwhCCv29TkcVKiFOpVejCn3HLp5+sMuSlv2xU
ZBsH/MF0V++QMdvBl1zU8XO6VMAkVJ3sNm56ycFa48POWbWVQCVub4oEfhD38RbrGG0sLHuzSH6L
LTLGtjJJS3KRH1kNDVCyaHHUSWJIApQUBswzuZeVnBxpe+vS664bgDx8o2lz537u8aBj/kHTq9DE
8HftrO3PapwWvsCh4SjQHm5I3+NM0T25n2yxfJMUijwzuc+jf7g3td4910R66JmfCidSNS37EEVE
cEElb5tBfmFmZsbYVqx5vSuiz4lbK2emQ9dZ7xZtbKQFvN48F2LfxFX1Qflo1BMibK7DL/JaKvSu
Hq7fMwd5B8V/RDlvZcOIAQKbZtSni8lLA0muEe7H7JrQvOOqEpQRO+KiPzyvLeTJnPV0Z2QUGfDN
rDnFzACd0sWBuZemHu80KFUCSJb2lqemRu/NAUBBF5VcqFtRzcwkcR3hqWNlpf530v8u96x0BT5C
AwxD6uheU3bfiL1OKEPRVolWV+WG8yYLuyh+LAKyaez9XSgTvuP9pLNIojYAyMV+2ywyBaPm2VCR
K6/9MOXNWCkRdEvyxTVz8TewNjJqAzcQMcxqJID+Pk0ANDgxnSIcFYSSOq8Pb4UpY5+YNU4vi6g+
xGXmsyaKZKPaYbfdZgy9YGBXVUyewZ31ge7vNBCRlMRAzecsYdp8TVGoaX4vbX5Y5O93tN9v/Wlv
IgogTtuU5BcEdsJgmJs4egoDoHCOL8RYSeU7X42t8/bnFrvgKRRK1gTAswrjUMgmp6fZw910Mt6i
1Xqq187Oz8qqtPj/SS/IrvF6z4ltyk7DSEmfcJ9HAQ0E/yBs74F3jFr065pr3IPPSIDAB472n8kV
xawcJ49oa+9PvkDvwHfE3lG84CaKJ4ynGarOkRKRJ9NMBq+Ixw7vdQh+1AgT7v2ieV4fqss6sVgN
EUz65sYGkcEejQV3wAw/cERcdxE8JgoYVw2JPG3P0y6lEajOBmo+pql0/cTtifXu1Dwd5X1560da
x1++VQEuXkau6PU35GG43ZO/k1dwwT5ccmKE3UL9UFrnsMSVEtWcfPGx5Ti3RIbCeEZiZsl3dX4+
pXJAJmR02LYDpBx3/qXsaG2MISGdI9Xb52PGeK4cCtsWl1tgCIWkCfB0xqOKkjZsokRGLyrZsWLV
gm3IK91W3j7blYKRzS/sB3M1rsbRdrI15BcEc/m5bbag+2eYx3ecl9swXkcFNT2lppDof26JOb5n
dAC/IW+aa2/oCf1wPfvlue6YjHgOAF64RtXQICAdv/vyFdfG7LoEBBK/SD4LKa3C8Hz8k4zbxjwi
jBqFV1uzEKEz3z/qHaBwbr5f1H2ktLdi+58uhmdYH512lAEPe2F3WfiYSos5kVPGaGSq4kME+Q0l
hVQTrpM9nqksPzTNQWbLo09iiB/NiI5M3c2KmRYpy5VcilIHBvExfdg+4YMuJXfGTbgm13j79cFT
sBC284qYeywd7jjx32CYt3e9jR4Rn8aaGj/B7HGMg4QABs6illG/lJ72IL9xxyHQ7kpgI//zP3WV
6ExG6AVDnujyL5amxhSdZHm0RcPyw/Qx3BMI1RZxjZk/WNmtyOsDh0a7xEkCqsApfeapvDiwOU80
G4UPgz9TttPlAyHX/WuqEZfzrbfN1yz9muttUiYc9k8jTDmTAhOvRGdL786+qxYiKUng67Ax3ojY
UTqliOlxJ6C1oRCwD3eQtAdZI2Sf6XvKQ+xBIx2/IOT0ukN1PQZF363ZbiKKuURXh1I3mgeY2eI6
ambnaC3sRSYwSM1rUHeCXv2uX5mNHCucL+xtvMZtGdWNK9cjlrXxLNDrzflBNEwUQQ7KpQL/jckz
It5ltDnGdOjoWOptNqS5XaPhgxEYlzKWF6iX2B9QJcTxArHlD4hajqMx5jMSjLryH6J1k/TKj2Eo
WlpXhQvL2hmiQo2rW6peGhQhMz/aLf1AqfYbIdLctaVd6db6Am2zMDqD5pEzDKT6cNPKTSSQz3f/
AfPkS/pSduJSclbs2PEV6JsNHTYHX//1f4F2jrj2XXR4mFuH6wd2jQYZb+mj66hTS2Sdc4jqMiqP
TitpdXSRfkVZO0OUPTKx4TzyV+zqvfvlrg+z9BB0mRsFj1eqePUKgFN4Qr+TQWXmRgEFvZtMnfoV
w6cR+rydy7M/uEIyiJ15XdUebF+4YK2nrjrQffLVxFdt9LRYe6c9EidZkfKAk2/1elKHo2xLGTMu
Sgxd0yvSePj4XLJY+BCk09Xgb7olHqofqBqfTDHfIUGLEJdVaAglz+NzHMWJuySpgCGZaHQ7cDU/
nrZripGDe3Dlb6krJ36lQLFYvyFQkYssanO27Aa7e46v6ZZ39x+/vsdh9fMoFrM5yJa10UCX6Ykj
WI7n+Bw2kzw7PISjFpnOwE4vTsXBrF6VobPpeS2t/Z0I0Eb1YSswKkqLB7dbZq+mzVKDJAVE4vXb
HOzZLuzc1Wdlu32G9ndHWxnwH6jG/sbmIEgwr6t4XaFRzAwqiYN6hqpUa+owWzsw/HhTpLgLVFXq
9WMoksmsIH9c7cLote9kJVK3KdW4Aa2tn9KqeNYrGc+e3bMR1rD2RrLLskKz4DbIxcvrwxg5//Ai
abVvN8SCINPlKBKUeIqOM1l5EDRnkDPZg5eoXaNXGYVDJybvVaAmaxP00to7kQNqh+7sK3+TmWD1
Y3ZpWM8EQo6BrHBMM0uYVNmbM+sHLsyeqdmCkjLcuEfDizun+t79rFH56Yx+uTtC38uBI3MUjXGi
OOgtYkVZ2pHABQ5Ajfh5oti4NvSNEX5zwz8NWH5PwvkXAcfGbFBVktRA/n/ymOosfrTo569XvvTq
FyJCywpg0KIPYg66MeXXxuZYrLwsUxYAGaED0UZbGuehocJ7wzA+QLVDmLQWm7o92w6F2sTiDG2P
l1Y/oINN638d4cxFTtIEFVrlL9jef6RoUu2f5aIXnLCPhytT17XUAM1mejNfcOxkmQ6cMdIKB0iP
6A9BcjKaNyC+ByYgQJww9YtjaqAjUtTMp/iEpxdauDLbjlQ6hwgTfUmGjLmAWt/6oiUMIHy7qz+a
CP0rvuiQc8ec3MbgpAEPjRvOh5YXO0AEGX+jis5LKN3fXjANn+J3T4bcF402hDk5xiOiQBe4tpWh
wJGCPC5L7mmytaNlBYbe2YnuAJWvstHmd+VuXq6JHp2NfwXOaoDLn5jhHRWQyzRYnhw1PPekRAqy
PwlrsJc8jtzx6ALToDaLzYbjHA2+6JynjOnibbSdFEHWDoREc3deBCi7hKAMGJ+/4Ev6aEgIkvId
RjQ6xJ07SjrHzZdBJ1rJg13qCocCEuEq3qcbbwve6uizwWE9sdzMIdqsr4AFCMT+kFltG0fPO1og
TSWCuQAk0mdozmpGfOVoGWFDixuP+MUeyMzHXeB6mS2lHGrWkixMd+TEafp80maBIYdO4fukVG1W
TUIDfdFW0ch4gaIArucoJFPpzy2tH/UnZc9k7aE7zTgTNpqJaiBaYSIiPXWc2jsIXr9aiQIyXZw6
25jTFcpglHnoYcT+vjEFGAggST7pCJysMjg8SvDBqxGt8J2OpMaRcJqGueo2ERrAgmZ2RZXS7+HJ
Ig2Hltn5DN3RfznqzJAr4gDRylZfmY5iis4RCoMgIZJcoe5ejV2zO79mi3mi4P7uShy3s3mOVOZd
TypxNUgT+jGS7+/CoENomnUTGwA74MzqwS/4qOaSoj02j/BpLHM9qwl2eHc8P0VsyQez5+3WcAwj
8jYk9B11bEXKhNKK+Q6A/D8vLnA4XiwlSCe4MV4tAUiYCvSVwmZCq/X98E/c3YVgNy+gJ/wWOedQ
PC+zSJ05ogymhR0lEIskRECNFix1vpc8GvL7OMdTb/8UGxylq6Ube6WHWmw7sZx2I7INjhvq3Ikd
tNejraWr0HTcY5eGyHoVSig9uQOs/5RZw1UAtuSqA8LIppmuYKfDFa17ZHqdGmwfKNWiwNx9Qpj9
CeAqzJtW0bEqtsRSPb3oGEmBtm9eVa/sp4KRvhiQWUi0ynuXda2Oic6XRIbiCJuc0zgPVuNomviK
ycAFAV8Ub00Vc6ezg/CAPldtPr4R8bdCuWeveW4cpMjWklik+jA/p07DoXla2mYx2uJzUyo8fe/n
AOcLF1FdNEaU/0XXjSYAVlxXY30C9tBoPsdRSIVV7O/5j9Zj5hXE6i2DdKk7zFy1tfabP8OX7h+x
b1P0vEVwM/Ga4hcApTzK6/qb+tnlflm5JQQNkG+JinIQ5+5twXjy3VHuvu5Rk+qnsNTaeU/83gBa
4jN8+deyAelx1azIRZJy6I6/OtaL2EYZqK+JHvGTZfz9XHDeYwoH2B8/2yv2OmA6brDBmRQLAO8U
6a4e6eeDel/7AzJvjQNico6rl0PtYnCFckUXG2CI0G9SVM7o+mr7v0RXCq9BT3UgBvYeOR5e7dIv
uouJHwHEPr/NCUTa02ZQqr/M2MMqVa1dtqMxi2FSjDovwzedogn6mfze3gLV0q+nPp+2H9atUVkv
BCF1Pt2UBXFX6sloWUfpjbck25KzAd2hXY4mtgfLzLTwREsB8uIlooYmkMj9p9bg9f1NfmUxC7vK
Gh47XRM0WbfMlLP/gVotTJKgoc5M3B4S9QEROFe4Pz5curkH+sRZM3726NqOwZSYkTIuWdVarrDu
EAdivKgit3YaDewupJUSOwVVrFEQUWw6Zw3d4aw8Pwqi85yr8oWNH2Yuuza7tFBR7QO4e3Jkm/Cn
dd3Lscs8sUS+ACw4BF+LLYN+wDkZ37X24KIJGiUX42fNCaFqljJut2f0Hq0lY3tV4L5mxF8HbrDl
cma1vASAb0kwdNoi6ICStfPTMCJWhQ4q61rOq6OocW+tS+b8d1O/VL7j27nUPBchEJ1Kf2E0bQdS
Q3SVsLFlqbIrJdtgDqPml1U6TJdXbuTiigO2y2SbhSLs245CJSeWt9GYM8RTo3rc3FsMK4bDO2Qh
dQDkbm2Gp7GN59F1GjZQiQhwiTGnlin4m5CJpVpx1uHnFzsi5gPRPN1F9Of+mMKh14zFYk9EhpnO
ct/Wp9whhCEGIruiye2SUpIeGCD9Gb7Me2SZV+exF1TJLqwFafMNGBzu0SlpmkJt2GUfH0So207G
fRPAU90ysAFAVEeP+1vBzUWZK0YTi+oLzA+8JZRGdQOSBZbbc4dH62qIFEt60LOoVhJ9WAW2uFoD
ixgZjK65t5Acd6xv1sfSVLqSZK7ptHpujRRMQggi1/uOkk9klPwyvIc2PnQ9aOm37BMFNDCDkO9C
LEm0rWl6ahqloE6Whowg5nAN5tWfilMHHCcWLRQOsvck62XDRU8P4cwRA1KHebMqxCKapWX89728
3TO1ur2wAux/IioYne0HFXstbBA3zVqHF2gFpbt2eDggKusf8cN2/CqAKWcgZGLzt5edZtiuAf7m
VlOu+69eoDcr3f5IGHCd1UG1xqf2MLChIslOqvXOS7X/jZdW46ccSB4XtTA7swIL8myQ4Y5xJO99
435gb9QEqNfY6z9GTNqkl2hfOgyjfauOrA6dlvBqCrF0ClvWTLfzin9AAbdpECZmm3JkxVaf5CTs
+gFrK6nmdHE957SiNbOpaB3Q4dXHtNhQidYH+Ul5mldz3kVxYmuM4kF+FGKfAPJYnWhwS9sHsCSJ
8Lk0qR60FHdHI6hfWXaaLrCz+i8cPsrPBj4SmkTnhlzgHpPISI7eXnSp7dfZ0nQ+ILplk1M67aym
Pq0ltapS5zR7456iJENRK6uPghGgvPh5ZfCs7/R6vFfHU/zbcspGLZ3vP379B5R8TLbS77jqQ1es
xDf19lrO9KMQLIpwRgVZ9FwILKioEfquR2klkzoW1oqSrX0/OLYKsdItq4+6AOkxH7uj3ziPH4Fr
EVpE7xaz0/F/VurWpNcFT/pDr1xsel37T4/7VDG+fcCbYG1/FuAjM9s8o7DELoBuk1LCPG0hgo2w
ozjQj1nygn+CDXbPFFMMxemBux9dUkGliJQ0AZSr7Q2mmHn7Y+dOR5eug/wZxeNcUgS+oGTpS7Rz
NJ1LUYLvuJW44tsrrLFlqgOafoOjOtK3159u+l5BqpyLKZYaIAq3o7Os7qyqpV30eglnyja3kV1O
Tv02CFD4GZB/DBU2Im81a9917oOTnq/BYkaHAnPOfSJNGx7LG02FJYtgDAne7xsooO9I3Xh0yM1W
F5PybIuzd7+9lmI+OeIFNr+VVdW9RGfN21d+4DP5bqnjbJsxCu04q47ecgEJ9ybnGyAdz0ZD0V3H
jXnL13Vv1Nhug6HEYV9U4CQJrxXLILjGflSilo5F8TuqTHRJ9e+U1SKxEKTyFugabZaQyUGqFtua
kGSA4SJb3nTkNb+HI+F6ic0R9kAs5ibn5RBl/yro86cWXwBkRoERRVOWwkbh1Xk7uAPayI5a1pvI
mV6MfvfB8FVrLrTlc322C17/rXOzZfSCDa5PUFWm88VMI1sVgF8d8/LQ/rB90H/kcIEBI56oAsWP
4ruaiKDjinn1QfzvmOLTOV27ZzdUCJFJWuqAr6tDdZQDBJvklc2R0KuCBDHtb9nafwWd3r2y8g98
MlJPaXge4/AnspY75tstHGhUds/ucWQwT87cDQKIktYzxLd9adIZxEDFcpKB/036TapKVc9ufpJ2
36uwYa0igi/ActSlUXaMQ8t1PHXXK7ZM8neew5JFhUMs5Pcm4gjMapQpjqSbMzUil7UCBgAfzyWK
P0osARqV8ZCAfgcqMzdLvJQzArWniIzzhRHyUrXftaTon0kuJxrQv/3HV1LLIGYD1ylG+d+gRwcw
UVZyoPWzrAiURIuSQbjHqikHGqlFyGuZFGt6itGH1D3gRx6ks44YqJUYNyWzmBnZClWB0J1N4qpl
suAG2by90N5IWrDFi8MflPT3xVbiaN55UdYJ93qnxlMdcpN5h16bKj7qjvJbHVTIxQDjGik2QeVh
g/Dp5DEzoBAUGy5kUr3aMaeH/qFQKgmhiWlhyd9JHHcD2nB0pndEA85urdlTfufZ4Wxmj5RcD5l7
6r7TgZEFqXoBrqLv5irnBT4c20hPRkUdTvzdWaSpkBZPe08A9/a8/B424RRmGjwaoLd3ENr2Einr
9SEQVubEDUgDU70ICGpeUsPZImKyThDlEjljoU3/tFbKGP1VgR35+0bBDxWqXi3CaR3JHXz0BjnE
9E+IGatLGbjXovKU2YolDrNDYOSoUwCe81nv9Tln1FEIVHw5/Zj6ZlQiDNfHJkk76lv0BCO4U34h
BIGlqP9SaZdnTx/a76i2YOHIE1+RTjRljSKMWj1+tS0hkHJXU+uN0gmXv9D7OOdb1nXgfR5D7WY+
iVX/V6BSp1vV54bMYhkxPLM+SMM08HkXS+2liMB6U2J9qaSHpRFxEe7SJvioJKoY5ol/8ZOwWWru
OWnqsccAitM72KZNY/LVJGSeeFwbaxNfrZtXxEk0VSjMnkM+oQUT3otWcExm2bNFNs2e1prtQz9E
zoMjrgCVkgwUWforK3P1YqRiq1XLuRAaju3Ut+MAr9gBowXJ/+2axqb3UrK8PQiAULuFlb+1X4P2
XiFp8jvvO9cbVVD+/h/H7zG04JrmTuWJI5Zifz+aZmSW2mVmVfJGbI66ggYhrlWNS9Fxk3HiCsi/
T2rD4ti9Q/beQ5xxH4+YZRdlkm3prJeDRqoSo3j/W5jlai4GJ7BicAkjtHQvHzbvL9H6z2yrfDXE
qFZiQF1YTzH2c8Ee0UiMjndboj9nm+HuJxalRLxGv4TXXDxD3PIYv19N1QoxZF+ZOObyqlum/2Xu
Glu0psNqkn0BVFKMD5CcWg5nF1JNjIcKDInj2BgyoYthlo5Ezncy1n3jadVaYQI7qeE2fsSUJwn+
GNI/QWsNV1vg4uV+M024L/jsgX0ugts/GkEjAy0kONVIgTGd7zVjDPPGDmQkcF6h2YSKM7sk8zUl
LasJaW9fygNA3abfH2lm8M9BAHl04F9jmJtxJUOMp8bELQ/a04k5ZHhtRrp4Mo3FryVKwoo0Zmv9
TSG0TQKo9lJ0D5XG7s9+9Vcp+BegC8ioAx5I0+28rZLFcKPaTYbOe1TzUFDa7WOsu/VMj+MExrds
NHm6/hBQO/P2ZD9Q2rAiQEjnLvXRtyp2vz2YyKiPgHf7TnwAHEZO5fMs/eQfKvfJhtIKCnKkhYNh
KDbc4HcNWFUaId8pR0vOHxHZ2Bgf4v9h9xD+MJb98B8Cv1x6GkSnsyvbvub0v9nMfw3CUMStAQ+Q
QNNRH2d33HiAdER8+kBK3n8dzoohqKzTEfRaW4rr/KvsPB2xV6+sJGPLapOdqXizKogLGeTHd+m/
c1mz9A/XUt/HEQKVIRx2uurT6/Dh77y3IKjCK3t03+xm7+/EFI3UDgR+ZgAk1RZPir3JTnTmHh1o
uaqjGYusHjtazRPimpFmn/M04Iwa3wLG7uPOx3rdlloWFoDJHbszNyh/4gDj6Cl4h6gp6o9oYLC7
P4nUV/+TKxe4QWmYfVGVG9Flw4R26/qAlYOq0RRnTWR3cn8Z9DRlFC1hn0822zD8nirv6zB+PXlz
VKUot+eOcGnm9JiMHv5jU9XfFQ65Hf+p/YCGDgtBr3DUc0apfYb20CWSM5O/wnBc2E6rFTtiROpH
lH/BD/ixTpsuGk8mF9PHkZ8GsBTNYqyGjBEfOts6cDaiobLqcgavdJ0jghmvU33bj9MHElaJzOnA
6BiLExHyS3c+SSKT2YRNI0jxhqG3wzCAw1wx5bCiqgqpnwR5S7Q7tyUpwi+dbqp0/XfoaOCkQYEQ
wWX6WAWQ3aKtalDbFlRoUB6IPtFuM9Ry6KdgmHeiyIMWEJomhSMh/cV4QP2Pb2BJnFia8zINVtOt
F+NByCoMHFpNZ41Rz68LO/plM1oYahqzCmdIHif0e5rjz3gnyBITCn6WqGe8zwmr3ONmTSelGgc0
b2OcCIdeEjIwEHGwEgyJ616STU7teCi83eoGjLu8GsSInoe4UJ6viBhFV0HPZ2XGVqS42UhXo6He
yPfkugVH4Eip+oBGNO2XLUBlL9j9slCNgAlwVn2n6Rv4zuCRkTnB+sHARz1fDHzgff4mb65t2oGc
D/7hLE1o6+AZz6I357EtF0FwIzLyJ1MeAgX426oY+hs8/3MtDJHSKN7kl5sKPWM6pXCiEvULVoC8
PTYIdBFD3LmC/6Br/vjv7aFhsn6OxEgJyinl7Qrd5FVQDnvVYPityNgqZkyuloZ4TUVWj1i3Me09
wYbHCH6pfe3gfSczQttkd46/i/m91e1SwiTAs3XajhXVl7DWoIfXAFtkYlsmAdzVRgnR6qMP9vBm
/BEXXvFQP/O87bFA6lfQLwpxZOMTMuUmT3q6AtY8YLklwN9PFaDKMV5WUUHs7n2egBtQYe8Ktr0n
alkfAqKFQUR5M4w388B0z4FyELZd6lzDtVKF5ff8PNawNNiMBsxUusd1xe8d/J8rdvAgFfvqE5rW
KGcnhOpi8ZIVCl9wa1Qs92kcgwJoXhQLzzWGH8jBbuRBQyRImsRXeYTvhkAhEKLyrM4e3TnEcPFe
4Q8hLGAT1dAdqHdWKO9daIfucB1PsPHD/O61bs8/iCK2YWHRfVwXO5SSzepX7MdpaSSxFIYKogfJ
JjgUjUXUobwcRE9TFpsgEDY4qFJU8TdAGKota2dILhwMqelrtmMbbsP9dGCDbtIZaU+qijr4pSRU
MJBjX314al76NZqrD7N5FXQQZ/GbbzV43pbY2MEwQWK2KN3jIRoItgutBjLHZAcORIrm0nmD4WsB
NGuWCaSxVv59lzGwuAIBLaaebGwKF0wRaUXad10+8kmCRmspY0qKvYCcrerGXqs7VgqOSN5TU+1G
yG+H5mk6zGy25SIHlJdOSO2+NrWTt4hwD+VG8VZz4Cyolj9rl++U/bbIU335EOIlnEzFaGrRRgIA
0UgdU885fdiZ74uGPPAbRyy/cKtBSZkOylfDE6tCqJthw2bETYnYrTBfeEKSvjfIibW4RtOSCfJZ
UaJHk3MmeFtxP6TmITet4qxXaptrp+OA7/iIPmiUsBz61c83zEaYrn67XI7IqnSOgjzdFQfXwsjw
lTjPBLHYUQl/Rh+PnIQxoiFJ+qLDzdJ+JpUIpKtB+PCFUGgliBMrmsu0nZlKAD0fD2yhYTp/q4zI
C2OUegs+0lKypk/Tsc85lbnkJvVCC0CHdsi0KM9NSTtD3zHQdGEivIN9xBZaBkWLNB4ccKTqW9py
67HbyJvyqFh543JH6lMVb9vOg8/1077pJKqZM+zzfXaUnXkKeURiEDqomIbL6cRoySz+k5cldpOq
tEDxWCP8RSwd50anWMcNISrl7EpH9UzFSVTicggHxItVUqg8qtNgEdlpoPPIObq56nUT2LrZJ+uz
mB15TUqdx9uEVkidzZLiOgdcmBNuFJOHKzlnCdN4JpSA0Zmox/tBphTaVhZVuJkkDH8sPVTkuvxD
NbNq8TGePpAsJfAabilU/44OKFaOzpPZ89QKtI9DjJxEnG/ZsVtU8yTzgHpIkmIdlfx1MBzgk4DC
+vFfmmG3WDcfBU46e+AsZ1o8Ba/7OTb45G1uEWXn+vZoSV1yZ3rUkqTv6IhIHwJ7j9MYZflGuTPi
2H8Wyj7t2Vsk5u8Jhn+uVBwbtrj/apGfZIeB2AzYpKLx4lBH0+jL8AE3e/RCkNbgD8Z6IWmWGvwk
49SCugwN/XvBkYH4f9pBQZMYuYA9r+6BZP++kmSIm0cSha2UcAlNI6UrZTzE/kuq2IlqgCxLBGw8
AsekyF71vMp/ctktLvJWzbQ2mrDr5sVPaRUwIe2Gp+FMA6MGoKo7ThJh70p5mX71n3CBbyZWc6Fl
GgYnbgMmRTxjvgyB/kzKjaAxahZF4PZ5e1uJzGyIpMhiSeejxpq6RUYSaqp4PBGTTGo2fo+r7NbE
Ves+tVU7dwoFops7ksD6MPbtadSbH0STEPYJ3ax0L1mexsEGRrvXb/rnXm7/Q5Yx99I/nVaWwY3m
Dx5fgJjQzxUF5NI08BwLYnoNJMXL78OjIeFT2h+bVvYtrenFWR+5i2em0IdK46WWQ7XOwAvatzA4
K0rVteBIf042duN+bLfenotu/nat9hGlEUtg2jd+4QUWw43BWTbzIjX8YueTdRGPemwx+V7TSt9n
+hfRr159MUiS7R/HhlovSbq0vGzHBCZp417OVd0AU8AhGWVnuCRKsfjRPXIw/uhrG9kUvUbIFldF
p/sS8ENzXpFRivpVn+qOOUPu1S2xGvdew/hMz10HtyS6F7pmpyW/bLjXojqeNhgR1upC2jZi2BBR
7TgRY2XoHbfFpsFnrKw64TT4zWS8/BgODytVdvymh+ZkFSM8Kw9ZoYNmSsJMjbtfUlcvdAEfwouJ
AvoOIkEdP0qSrDn4jWdGAETfMU9xDz6mgPtOaKXMhOZIZkyzqTMjUYQFOIoRxwhhhu0cSptDHHF+
81fX4VigjgSqRvVuGK8kn3hYLN6Zg8Ysc48vZya82sdvtU/W6RhSet5d4S89kVcT8J58SKxbvXG+
8dllbYXa/owVq0Os8OycnJt2MOjYEKBKMzCtDFxM7ouNIZjccTQ3OXkE1AAS3HrUBABEclW8AxcK
mQNFAATGZquwH6q6kIIC934sK7LW8UI8q3BM+Oap5pI6ebzskYPc4eMNSl2XwX44O0aKHGwUWfaM
IspXd/8dkqYCDWQWI0Y697XahILU5lOmPwtC9eKLKc2C0xTA4P83vhXi1E3iFpuWufZzarmeFlG8
SU3OpSZpYs7GNoyITYOunMxHUNBFYOBH0PuwUigHovtApSCNeWPBxhmg920ELAs09cHFfCLymA0X
hO6jGOvj7hLmyuiUpkr/u7v9BxooBDw4+jBLaQNJKH+m7Dlpehyliz3si1NJUIwuwTxLZbi1EepS
K5Ej+mIvHYUZD3CQS3XEKqWBHVkybgyXJvpbuia6//ckp/58Da3YxTu+dQjMaoVhylj+VbXjivfc
8ErniMW/MsgTyN0JlFt04ask8AtctThTmkCMiXjbm7/cK65bztxZgk0TZTRQZWLAgv94R9kTYl4l
mI7jg9QafEJYq0oHCL/Vt4ijJsDrcomFcalv3wba+JB/BnAG4LVydk1h376na2vzZoP29ig8q/8S
/HRjPaOkHxTA+wyHCja4XQ2+x0J+Hf0QcjYug2sQTodj2hep9eu2qR446CzyH6MNBtXEF4nL8yOR
vNNGWhFiHVePiiiVs0R023/u/ZlKDHQUo9F/NrFFlSyAC0Hhe2XbB1PkwB3g7GA85jYKGOF+3k2H
Ei7/Mm6yzVjeEzhYmtUhUC0sbY3QsQFgl5au4WZdpvyha2CKw1n0rZ2EJCd6B4t7x0cLLJNAxz15
NKIm+fF2cBdrU0SrbQAGMefbe/qzo0y3ZuLeXajS2JyvxoxHeomoC5+Bw28I9WWXuLKTWMpMn7in
BymsvcYeisCSOnJSWISZBvs5k0zG9T3XYp+2VKNMMN2RrBVRkPkbtv+1aUJw8rIaOYoCDDgd/PC6
1A4vy4SXverdIfuL7WRZlNIsmV5vJROnBi1vAhaU2tSqKRgVEOA4qHvUf88+Rsd0A1Nc6AX5bvjP
BqTJQ2QmgYXpWjI8CZS4w264H9Oleu8z2bckEV7jtWbRV7k/6cmLN1+uuPCzf6OIDUULFJW5HoW0
QIk8n8fSn3WzABkcR/73orqnO3LHp8GmxkOmWzZamDj7qy8WM/wgnpQ5LGqY+nqIFcANjg/+H2rC
tEEPMgS/ZvNxKMmWyhIQHn7NHjNNdJNtJk7OB3AEupiegasP3pD9fymAqenXniw/5y2arG8bUVHv
It+VYY++JMgP0CxyloIXiLAqcfCA8jrV6Qcy3EwU1Q5NEox9HHSfxgxmhpG9YW3Rj3O7ppF2C6Ko
J+I3zXlnn8wQXjLWhkBd2lVkiZL7/m1dFcyhmWVnaE0reM8LAEB/H62+tywMHr3k/pIHc3YTdzIq
UC/l/iI3iDWaL3xmuVx5V44TEgBCjPO1jM6NltgGIkEZmCgkKwiH2qXJkvdIE5X/TpHquQORrvHv
51TJBoktxdCkDMiI8MzHlBDPBDFEY4wEuqlIp6WZKbGNFQOJ9bdiq1byDgtcYBpyLrxJXsdBW5AU
oiDGfkMnXWR8ibNmEP/c3Osb70zAiD0Yl74ZqKOHZu5FxjUZIDT/NRa1tzIrvejQSpufrd+Z9ssd
cLWBTL0n+uQQrqzfnnwPcuaDkwohY6fOa9Ies0auqVLlCqPWrqH98hh4RgHLcM+ZM9tPlyl3TWv4
4ExebCi3m2HiALHUXOk+nDGTb2bzTGuYKty++Btgw3oy4sRpx645KvNysIpsowz1V2Xg3wZiYHlD
u1DIvl7CetVIslPZyVGDPKbi7QbqvMWVwyi5BnpueqDnJ91dbDOiz4Uo3PspjclRckgMPuhEztAd
fDD3TooltAgJNGqDtCkNbVDMJYh41Zrye3VDG9ymzLwhveGzr20WqM8ThAXmUvCZbzYwtzp/CTDe
/DGuW9fBuXGxKdEnGbxs0xhfQHS3WztZBtZH9YxYdgOybkASbPJoadl80KUzwSJOaPS1CAlZHYA7
P5/aMNHX/Xoye9PXc64sN9hEiquE3oPg7KF7jWaGHl7S/akAlh6Y2QIbsVFjy2SSNOzn7FDwz2gC
eR/QV+XHjSxe6PEbEHRf77091VPD4/og4G3KvdKORNvksTNrU5p+7nk4ZW2ueb2MY97Oqm34vuwl
xV3zeLvCho0U3g2jTATrQt4lxwReX2QhVAVgt/gE6aJeImAsc8RUlxDw6Jh+VQ7VLTQo1QMor7Jg
FNnv75HuD3/OrTBfCk0bynaTcDHtzjNkCMpcbdYsICzWBOQFbExSgR/ywbM9XtxHb8jyTX5yTCz5
9+UZx3T8Obddgxg13fAuvcc9vaT5Wv6DENwU2kI6cMsUE09+DcrGs0qaOEvH9I7z/9+EcPRJisVi
S7kQjV/nOhKLWvfLuHFv2ZK02gunlsz8EVh5VEVCqSRGaQLJHBHuzKSjImE1lYZIPg+ABn2BMM5b
5Y2wGY0IrTrPDXe23kgTy9aCnXV6LAMehuEo93bS15pBTBgK9XnhP7G5oJVjro8mur8TzPz+yBTa
l1eWEIBvLJcpG86Z1vq3FUnTaQ7iS+OsGTwUcwFK0pDDJDhhyLZXXiAGdxDmaVgMfS4otupRYI4+
+E17hz7QY7RZHcX2ums+78fUibS5CbhMeODeUpUlFew2+CDTbk9kkiZTvahFiN4Gg1WsSZrlb2rb
/htiFfemmfQ3oZb0nPtzByG78L5tdEfCwhY0B8dQXeuxhAIwI9pQsfxwXWYFXihrFv5WPXTbGWM1
pYkVxF4bFln4RMgp6K8/lhsOA3ds8TlNJUXOViu0JpbbVigi+FN4+ENyctvNQ6X4YjFFMSFhgtAO
P2Ywe02weEOf8KrdVM6pHYJ9mvA7oMLzILbk6tAp2HWwSMicO2iRtCGGA0M1AxhJ6Pm8uTbTqtkq
ZwwxpzGJ24grUo/2c0MrWIN62dmiprhb1yU2qOp4EfteWQqW/UlE4TYNDC4Gg2zPOqJYW4APGehc
fatanM5oS2/XrxpX/sMi3LCLZsVt65aCk7Lxra170RnYOaCdYurtk8KigPmCAaFf6jggoe6VeJ3q
tQ2cDpdtrMg9ABDRj+86yApwBRjpJ+5HySw4T902YyQ43iXlqqK6V6d9gnRUQCvfiEIlC/UCEM8p
DNUVhy8rmgf1OItV4KVZ1aMmIXmwUg4JmyLZ2UONC7Xfked5ybial8Qc1B8B/qbhF36mgEAsaMEi
5Oon1Jb3/mv/yV515ljUh+lTCkK1eDOhQOR9tyTyXuaxeXicRe3/U14FVCw9QEvJN7I305cHc3+L
HajQsXsv9V2kq4Qw396NvSqeW1/UtNHewZBXDSWJpM9WMuWtf2OFAwzgCXaAhyjAzgnfo0k6xOkp
e3j5ZkG5AcNpxhmufT7FAUf9YdhLoWq0oAcbfk95LVAr9DU1tnc+N5P9wVUT+JQlFJ8a0YxyjYZG
bchwrNucXc9fZTi5jr5iv0VWWO2gEgrNoEd/PtVL2oWjySreayX73uMZrT1ScHag07PfAJWuE/T9
5VS4NY4E4kujXjqt0XUHZ8AEqvMTDEzxFQQfDQYybpf2v2sMgPyF4tpgxuGTQ7JTMrej9gJcTyDK
EzS8320qvA/bQNZsItDlO6l6DTuKiDennEwtCY5VFiDlNcdB3ECe7+dOFE1usyMu9g3Vrrl+MuHN
bol/sOKxlJ/0QGlKPOsfB5oY7VdyH089qkcGZhZkpZWbS+q6y1WfhWg2ukSOURFMiD9V04idCozX
1U+W2Rflk+B+JHMbUmHQCLMPLeYlKM4tPM3drpSn1BgGjxIJACmM4UTaVD5v5VQ6CP3+svBdH3ou
RBVg4sgQAJ9m17uwIJ8+lYJbplYkpEN/7nskBg/NA8xxl7ek9Dp1wo+grkVytWJCyoWDO+blEopp
OKUj+txCBPKKX4FNONZIufmtGPxFMhFE15f3bxVqQgtnj7qaDBdrIxZUL2jZ9qm3HHcYHtrSM2dg
2kL1jEAbAqxcQIbdeTuQ8+jh4rtssrGn7IvBXckmeA0eiQIazBeqV0CVEXXM4BfRdnVjQ0bT2WqZ
kbT65j1y08pgHSyxxlmpgzLQJC2E4ueY6jSkuxKRQForLkReKooBovIrB/qv9+j1NwmGU4XpENbv
hVQRi7stvuqM0Ii2fcPdGmiBAFoGjDson/aVRBdD+lqfesmCuuU083UrZvjT9rMmVzB2MZBvcasu
+q3IDcAGtxfDBSICYHYI48z9zvV1BKJnsppvr0DYJjDXF3NEv4LXTTOOXHHkfiilJ06QUGq0ZxBK
N67rPIdI/GXCAEnvRGbp3ygeE0zhCrXvY2eqHqbvuTpdoRzAJqX9sGkF74fjr2PAjQ4Wk5D7EF7w
Yd/dv2Ftf0o+A6JPKX1XeZvIU+rHV+260DFiqsyQzF8w89gWUS+5Y2eq4uLPovjjY/uiZ2rOS/TZ
5dgcZ7PxWO2xKHHtsMFNIct3mpHN+xgC6iFpB4rN4izIxhUkgojjaNjNgiYEjXLv/+8K749ZHEmI
r14oRL/cLoN3KYqlQh6VCPpzqiIXm2d813J6G4PW+fDTlwDPC/DU/eFUVyu+EskAKwkEOuRuX3pG
YreZ/NJ8/Bt9jHx1oP1LeaLj5btiFeF8dU2/MgNvsxYjhxfjv+Zw5Huf7BbppUuKOIzej3dt1UW4
YqAyq3Q9ickGKrz54OTpkqOIHYZCg+FWVVaE6L8dsbpf02On6okuoiSIoFNkKaxRzDUYcnyzVaBI
mYfYE2xUq4Ql0uwhcRh0xArJR2Rv4tzJJj8xvaUzBdl8D9V45rabt0h4r3ggsEYou8akKBdLiWnP
rwAtASJnTUmAgyxr5t3ZzR1FjNNHBUSwwEnHFkqlfwXHzWbMdsw7kFE0L1PzfdKNYSFEelFr7olG
A/S/WFEa9GsvZbM9hty+8yPVbdE4fqtj9e7+pWPF1NPpfaDFfhu3cFeOgPLF5pvf8TbiLfPPHW6E
u55ZdSNPpjQCvIAPVKmsPBhm0MSyXt/zygModzY4T595R47QsWF2DenjfELXszcv7NUYXUxGDEEw
F+CUDkddZ9Kciy2dJbKmRgrop/qNpwyp7JSP+YLAwk5wLQEZz2C2oPn869GykbPPqM3lg8YRoROX
VOBjPHXj5ot/40vCSmT5CTAhBYEVqEGp5R88s5/mdMikjDILRsndZGyroHNEaBuljkV8cGzsPi07
7JU6rwGJHWPjHtE4FkdalFBXGfAC01wNZKaZVEqVZ/6Okw678u5Htmvcrtce1D0hGtPTlpSk1YXW
HDwNuqKRF8RO4qwn0Tu+CXLd8xfRdHS8zwMdDCpX3QIdcaMPdyLPdT8sG1xHwfUXAAxz8WFzb0gX
H5aJOEKmGIwcr9YUjloflj5HXeX7vDEqxPj4L9AQyIpbLsKyx+17rqaaCtlqOFUjAuJQ1ytvBMph
zE45CqFIvFCMLV8lxxqWD+MsSNAHblc2BTVlYK83IGu40OghNDSx6d/5dpW0f+J9VyneMipO/wXU
d4rI76rzPRwq0pAwfiv1VdinhTjLkl+K/xij/N/zQvd4u8ix66q3oL5xV7zSFmPPJek/fR/6LZwY
2ir6jPxVcarUWFtcz9517c5X7w40M+R/maq7LTUmIwApWLSUuzBjonWOvqzR+PYBmPfvGvelbyqR
AY8QHb2lkulc96aikomLHH89g7lrbil1F/+ckiJhX2KgkcZiStI4fN03Mf8aS5xvIWyEUFtm7r7J
4xP+1iR2wEuQ+r6meoHH28ZWbZYTzMfS7Ii8AxCSOAfn9eebwmL/ps5Un/5dWySdO178ycPtEDJE
8gHncU6KLaKvTgSziR8XwvWzNq9SUf21NGa7yajcC8+q6w9cOxoIMzI3iTcUvXZc0KG+/glUuqbu
lHD36N1D1O0/KQiUpUFkhGvratCb8bwMwnW7H2kbSP0d/kNPaDMYWO67etkiqlt+tQZnueWh4goq
81paSWK+rvy/i8jCIQmDHjC+bKfOA2brPSeXK5e3Fycs9O5uGs8rHZ5a19CZNmgjrAeXywcQhqah
15IXKm/SLrwFimzqyMJpGEXQRwUKwa/iGzY98r8pmyIW+5HPpgyBqYbhi6SuGlw3uEbIYVzJOlZ7
BFhjxgnkZle1c2O8kXPDLYmSerfXaqz4pUFMkg6I+NULh2secIbUuD8qfxP5YpDDKcgeY79vk1l9
t5tF2hJsTtnPfX1j+CKlPa4CDeNShDW5P8J/oUBLy7i77b6C5/OGNxsIgtYEUOKmBVwCnDNFoNZH
e9yChDQXlgjg1buW1md9I/p6VZATMOH1AR0GxutbJtoCByf/JaeDK6UBpWsJiQ6+93qPXAhDsIeR
anfuT3oaxas29ql7NLvDIxUb4GvrnfrfzCGtHGpcwAYo+vyi7xiUN42U/Ak7EcThU5YW5Ahiu7X/
n5Z6zLAmKUHpdnqR+BjjG3iRNz1iRufHWWpB44dsTgfB+Hy/Vv5CJPpLcGR2ANPwJKSwARNIMWp9
0T5wF0eYWFFhiVs7S29mPPtm1pIJZKS1Yzugn1+k2NpGYO6ipJtx7cYiAGNi+BZtRiYYNS+ev4Ua
xp/v5n87bFd6GmSV0LJgb5l6BBZj3H9Uh79jlnsdOYn4HGpO+7auo4U5OrYnEogdkgMbv+tAlr8s
CLHkp6SawX4bHMENPC4fSQsWPOvn1BE/m2L0C9Z63MVpKByynlW70CfwlY7nDx1f2s116lcgLDOs
dbNFtRcWIWHHy2SPomaFmRerj2k/w51/yC9cJ5uBXWlLloO6Y6gWMn5AUaOl5InHklVK10QLULWx
Ix6hOIK9Wf5aBXFKmxL6H/AzMphKBpG1WQOkNzpkVavpYP0xGTEGJDXGdoMV92FXjtvamga6/+Tu
0/2xWOrVS6g0bnE5fzctNTfjy2WsNDqgCqzMuuwZfmySEXP56pTZMK0aj3k4b6ZhXu+YooKeZlhW
eW8x2LudIUtfVodNjC1TgC+uBa5TVZe130ynUY5HDHmRMXBKHmBZAoWP9t5UsVHq3ZaFpMb5N0/e
w3cf4n2yARJYO243E40+MvgNuqhJHsYG1gXpkBd9IN6tMdMNEHEzd0cogPy/qUCJgfF7wn3XTuVV
H9fSk8TKunmXirqw8ayI1FT0Hgzdk4Mg90pJoEdIq15ZsGwfa0FS7N6lzgXjkK+ZB6/m4l9qvvrc
PQPJuxrLYUy5wmYAb/GV2IQO29VYeNZbuhjFCh8zl+k40F9FodiJT93DgY0MH67U+5dyi8/Ci7ae
6YW69Q7rqPvaIuFjvRgWnNoRBfez0O28NVhdDbx+47swKs2iJ4BPP8u67hFnHlfbk3815H4nN5VE
YidrGSXU2xNgwwwdQs7BKbADIzmifPzJ4xSNBHL8GG6wYlBgcXnqwBXWFhkxyiR20xST5ZKRF848
JsQimc5taIVRqqalLGJRw9uxF6uSmpzahtItMxHdt/0nor8XSmJ3kfF4iSgg5hAg2JrW3b9m9exS
tYDiZuKXfS4qQs95hORhRc9kky1NnM8vxO+Vk7kQOKfTQqCV/qgXTvJ2CEkelj8oqvUJg2cZoDM2
NJ6w0vb7nirT65jFSdtdm6pfnG1AxosWoyJxrOmzUn5UquMYMctwIDS0beQzAyCzgmQ4m4YsNPme
ldKlyiOVWTkdV+Jnn7gYDSVkvEGgjBPJfkm9AnTyw3+t9h5+gajlPjPz+4RHuGPNaUXzpS/YFWsP
N//J2APICyYbtREPh+pZ7EO46bWvsIVA2fIlIv6Axsb1OnnEzAP9qzIC5wvYtfVM/i7+u+Neq+Nn
cqjzFX0+ydgrnSleyoWFKW9Q+vbe9bE4StGJfgmdH49w6I2uuTQcFtZ0ot2qkH88nHpwIR+T5rp/
gPeF8D5b+mMrSM8xsOCZ+DNMXRg1MobSdwbEOb5pvzvw70EtfHc0zkmdUEVyRR6lALgKf2V5Qd9k
mH1W043920thO072YEpW/BoSicBBQ8cNZeOBnf1a926lfPHu1YfC6H2S5FjY9SJsxEx79mglH/2R
fJSI8hyM0NDsSibM+9Y1AyLlCr11elJIB8g6J3yZ9g6HM2ILf1jDiWgfVSUFTuYsVmD4nOCeD1z/
4udRzuVKB1x9un/SMg9/jWupOFWsqGocI3zXRX91mwdCZqE1ThV/koIg1uCj3UAjEwFjnfND2XWg
ut11bIARlk0h4KLk9f9FmoAE2lE+J3OqnKPRxTQ4uQzMZeNGmzzSdV5pNWlPd6W7OQ1PKXTJp9tm
H4OoRSFAvm6RtKwFIfwJIQWwtHkHrdwY8CMwZj7nu4PMApSe42B2nOuHaYjiSw2GzATPgiDkcmFE
0ROSsWtIL0KwNMyzPlWTJoTt85JA2MSmieoYGxUaF8+VuLLJnOZS6rLzcFFKEE9peqI7g6+Kv00B
LVbh0GHqCwf/dEmREIj8tDf1JGdFInQhZRWIm6lJsPh0gP8DzcTC97RE+mY4pxlac8+cqTn70LEQ
bIjfGXk/rnPP819lG6wjXX/eTf4dP2DFpGghkgCEcpNc724G9iHG351FF2C8zztcZZpdO+L/CGTT
snafTbJnFvIB+iKkz7GjXCvbyAq4FRIDceBYvx4Q/YnCvkN+FeOwfyfl0JLpt3PmHe6M7GdwBMHI
Bp2lbg5uLAMu+v8wl6vpUDNv+GeQv6uECrCAsYJ8MF9CY3L1BMKPS7+smflW9rRAWTtdVBUEbAws
csJuxG6DqBPLOgSWJ4Y1kB8rNmZUkcFPrXCWeA+5aktB8800NrWjy5SshxWXxz7Htr9HkQ/RPr3E
p4tqUJDp8d9P125dMrOkRc7HpubM8UawgAlVdwu+l3JP8aI9A0ekQpflz3Prix8Zf691jh4kaB6Z
8Twd6chwphcepWth2toJWn41mdZKjDCDKur7bKyBFkFl4p4mqp9a1YfarlFFc8Gqp0yqdfCfqHxa
kJkC/mza5eIKLVGkv2oUaxmIlBjZ7TrQTP2hEqArjJxVhvgsyWftBnXzUX93g4d/+tFLWpyAF8ee
R8UZqbKmnFOdA4y++9d5wmJVXZJCH51Ifb80wnZggZZFKP75p/t+TpZoivRFxdA2duj9urWZDPoN
yLu2F44s3UTl7Lvtzppxy+37xEBWXBsRZ/RBDWzEZntWYa+/TKUaccBsYOh4IW8ioiBzc6YLhuLs
wsHZOyfaJ0UxbD5oBaa+l4D+H8gHG0zoONHMXdnM9JPX08oH4KMRQ2lYrcy0hj6A3zL6CioyUJxe
Jy0BkYl7FAgKPayikSqYr2DirGldTm5Rw9Mc5M7usufHpJ7EaQZ9QAOBemVqv4lerw2j9zid8vnj
9ACL7UGOwr5QMJ+vhthETYCuIEyshfpfksMX1wzIqrQIvsdEkjMUfNi+LEaOCfTEIBfLfSPUczua
DjsgdJFt6reDpKQZ6GTLSWiw6jo9SAIX9p7+w/RW4YAK8hYpfZZXwStKfvKPFExiLOMNdavPGexA
9vZgHlXm/CeCsaWew0xwCQmLs57np3n09Y83v9jh8rFhW6mppx25YsvSl+lENsOzAjS/eC3YEKSB
2SeBFFNExxLucb/ty7xxXy0ulgx/74Lzp3PJVqa0OdgXwaWUHh/nMGrTR2EGtLK63KEzjq5emeVe
2Awxtl58YXC+CFXh/el7JgUzW/64qwaJLtdDH5I+VwJtHGYDRKW9sGlgX84YZb0+60f3jYOwXNOF
gmBil3Himlh8sl5oeSxuNIw4lyrdfh+g+cZdyurLvsoUMrOXy3i0Jhse7AtGpANonl82QmH898+v
pjTSkLWgPVhQ28L+lpEqTM26drlD8zF/UPRyNUSioq0eTgWsje6+yCLp4arPROnHw7i/BZnCYdjL
kdMEa2tAFZetSTax00XkIXihx5GLjUrlTNrYavC3J+p8EmhLmuR1WD3PSkm0XAzB6ne+zgty+ZF8
3phb55bqfZv+XOKEbxefg0EQcuBDWpEPiIdLCBWW09gIND3RjdisU2ddfYpYrQPY5p1quzqaDb/b
k8rConnssjrrbleQd7ksCvw7zZ7BUumef7rt80CMUHIN34bRLm7knJqyt9XJJw0mI3QBwpb+QYT6
DjXcLCTOaIsJke6/VD02JyY2QM9cW9/xFhyRyUijWA63QS4+31bVLo/Oia2pr6oyWytQSSaoYklr
KbRFWvAFxsmUNk1lQzm8Od4aQ40X47PFlSnGAPTVuueT1zUrb+5L+3Cd2ugUhS6CCdDuiu7jhdGy
I4pwIMfo7cDzIfUUm9KQGnlxAg+0qyNosB0p5s5C8mXdj5v1NvA+B9NypQ+GDLyFY2OYKQNo5vpE
KR7/+KNi0og4LDylDfxi7ly7FMWLkfILqP+qCP6N8B8r0KUyY3OyQyVkKVL4QDcFQyAyRU2SSuZv
GfyEIUD+8lhQbrFMT+QzvXpbpFy+x4gFNYKKsgVJPEDaQtmCGMeTpHmY+86I/fmZW4kyhO1zT9qD
G77jYNEwRAWmm8Ayuo9xAAZL8nt3vSnWBpUXq+fRt+Pa9rar3NPrrHJHPo2Ach1ff/GiThw+NCbx
NWQYIcv9WpyQmTmdqhAEK30C7+RFzDbdwrjDcvn4cBqBt1f/7prWYaMJB+UdnaniRceNWV/4Dm7f
xTeohsOgQ3bQu0iHHHGk1kAy0y4HL4LOXUdNXYYp7HEHl6Ap3AwzEqPzzAaGY7RxQq8HMTkfCi6y
zaa1wuF7wLDsRDI8WqbHln5GTzmeFv8Jiu64o7ROLrQpqdX7kQ47rBaIxRi0Q0+BhlYEVkk97+BZ
98IF0dKOVvx4qnBuAttAGs08UekqipeCxhJ0crtVIOU10y02YCyZDaaTlGP7zL2IbAkc//vnzWHv
A4kdGNrhraa3VWp11qh4VZfdvjqM72x93kDodb7z6xbiJx1pi6us72UNlWauX+0OjRpOj8QC1j5Z
ZXdjDZpNLDCj95dw55nYWItXwjhi0L20/uEBt/KKfBvrBAAvZSsEB6OL4S0Y3x+RN5facuKeioly
e0wi5XyRLYiC7mkgjVfKCL+SGARL8Vwwmskw7AF9KhUC6gV5GGJcFh57VGfioTps9f3Ji1xn4Tcg
isSoGPUMfaihoMT5njwisaEBjg7XZVeGIhIzhp6F8qxi4hnFU3/x9O4NssZEqZoFQiSuHlQHEkRV
OzIP+AmtpUuuS3BFH03o23Vi9EsDdzF1oKlM6HhpXpyKw6UUKAmSHCMkEMmQsdbdn42kU92CmdAW
o8jm1uGISVF8Q6u7oMWWu9za58GPMuj++sUDwenJuw2U8v1qKknkL3GJwQJ2EoYq3km2Xzp3n90Q
QQCt8/ihFlwVY3tr2bifqPbHbeqmIkBoRC7/17xo7E3aro9tev5oqRVEXcojSUmVoVMKXrP1RLoc
q9JFfbFxtHjUKa8VECe/q5OfVoj2H/kX1eJVet8UIG6d0FtIb33ZUwohfwdZ0aymJLmbwPkCnhdc
C0tYHdGPhOYOQ3CymuJnuffMrvFIArJRf1NtsYNObrfU/FbW8FdsibliecAAtSdBsSHUdiQ52W07
iOTM9QAACLYU2gRCCI6HnnQE5cK1mwRFJhTnHe8vIjsiaj4AclP7Uf71IUqgVgpkLXWvsdY8vAiy
q+f/lLAu4ZAzFAQiq2fMmQsCZDWYt1RuIK0rsx2vXUZHN+Xg3B0CUQGBNxS1vQQMJV3XsknrwFyB
UsVFFSkcGXWA9hlWGV4sLbKT/JJkyVfl7+/+D6Olxc07/eli3IkPiHg7ZHtOIiBY0qCkZrsBXKUE
gvqYv2+6qcg/1xmM85Q0Ux+IbzIvCZwRdycyMxXdjfEJY9nm5Hl4TZeG4d/rGgzqVBFUNcjEKjY4
qnljkhtXF8udr8I8UDkj8CWq/DE8ITIW3P0xVYJLe5ZFdhlQC98gQJ2Q5b07icYXWqejTXjjepqr
OUWoYtfnk2dLX3z9MtvX5Oh6N+K77XIzgAAMP3vD0otU+5uoQNusbWrQ+tZPaKuUt8B1dshqKJgm
b86NA/2hhoWNOYsUUj6O0uXvYB8dkRsnM0aBfHJ3x2lbp7VM0aOTU9cpJhgcHNY7k6b6ETA0dq/o
kXsnq3vCtAQGgpp2bfJeyjJpDbPxiLmb/chUTQVxA2Y/iP76styEL/dzxyjbXnmbCSaCohaLvZkC
iNK4+4N/xy6V82ua0ZoduXD0IBqhJgrlmpcMXhIUWD5ebUGzwyMlcMpXRpjGtv3fCbfGpkNKSMFn
QGw1/bDmQpyODRVfLlY9E7vHv581i5MIOIH/74YWiV6RrH0SOp5N8SBASnj4yBm8lLAx9syR3wZ4
tB2S95Ql1fyaeXrh1S4OJk3nXt29QUrO6S/xwZjvSpcJ7s3sk+lY6XyvftEYeFa6FhTrlTd+B3it
q67Fzbh6V5CB494wdtz6AVcQZVhsPGs5mOSTwgyt6Lq788tLiy44GFWuMXQ0AjWfXqozJEu+Hucn
LjFy9XHMG6WA4jB61SI0bUGmY5sx0SoUnxnKdhBIW8uOkAbZmCnedFK1v+WtJ16ScXDDnJhI6v/1
M+OJvuEgxC9oHHW/grVt63A03Kgo2/KLmEZ9VBKXO4SCywC7sFYrRmlIOARtt8ImjhLHSSw87eqC
iwZWFyGPN/jxtu1+ZZTPn7YY9Hr4XVTaDPbYKWnIGqfAGxbx+MgzGpYlv1qg97bEBo7DkYGDjPMb
QGfmWHj5wADNkyhXGvqUYsVefCs/IvySSesU/pyKJywHCzw2mlSQEJu8fqQr2keuAMIjDq50hv5+
8xC0g0fecV1pC+7s/ks3HvR32x0qDEEyPB4cqFRbTA8ug30R/cC7GR5zSTXXrtBqnvAbofFI3yRq
iY+SXvGrRh10iH/bI6y/LBGBUnwOY85pMhfwT+g+RF4rbLTimx+Fh3Bw6dL9LkNpK8ITkjN//GTC
MmQ4iQoOKe/Rv4zCHttqcVGLONDbivmuziqeeQh1vNoeo1LpHuoXRZ8Uafwl323RUOjrxakfQ4Hs
psHtpLqRahg1TiuTcD8gYgeq3dEKwgpAIbxUThwCfS/IHsg4AidSrgAInLaCDPrxXkhJSSNNgcOl
u8//QeG3M2gnCeiRjyX9UIgn46B02pl6kj1EnH2egjEFI5J5zCil+fjlQrjc+MloZQ7/e+7k1zuC
wU/N5PrDQJulv072rfdAspPhnduDvV1dkNQka5hpUDb81T1FNZD0t7rivdXZUk7qz4hM5H4Y6PTn
AXeR9klFEJGGgBA3cxL2yX6UXVUNcT4mF1b2PEZqhTXSeUkNBS5HPT7Kv0Jll/vw1kqzUjFhskSe
dNAP92st/7fsfDJ/aMs7QCmhUOo3MOlF46d0W/YWZQdLChwMxWK6DMNT+Iglz8nwrmjBPaJkNfN9
Y7dhjKO+Q62RaBqXYbd1vexRF5E3qWCGLGwbMXqdI8LPMH3yoL2uc4Nw23VocRcqkktfK/KpgfUN
lCOIREWy6gLDGZlNCXI0QhL4clE0SnG+EVYM2IkLtAUNM0Gj2aKDm3L6taRFgFR+Mc6ZntJwHEos
2vpuHWFigl0wj3wXKNTb+3xTr6UuSYd9706QMlAkGK2lJB+GIlLS7dtGUBBP72NI6yhujtVUHWQ5
SjxXlU03hHH+1oke87L6h2PcnADmY57rvK0YQWGGURy8hXhGFVz37TWLgqxv49CAb2M0RXjF3sIZ
OwNCWcTGN6nHbtkMFwg8/5p+0NUdGlglBuUA+UYGp+gv4F/Ep+ym0v3ku/xu2grV22oxFO+OKh1l
PBcHL101hDqbXid80StmxPZRyXpMrQI3LA9bMVqDQbz7GCElbaDTnr2M709pSeciadzMsRXpmOf+
+PxpAosRGQSoMQ6DBa8RM7Y5ELHNaiOmFxBKXdeiSpBFa3RP6CROLJZ1dEBsYUl8Uo4s07Pp0v6F
mUnE9zDSz3Qqwrpl0lBbJBJHpZjMWs0XWGp6hwCPMLpcinwJTh20I5um7w//Qj/1Ctc5OZSNwVcc
s8SPp/MsXbYSW23RPORyi1d0sMGOZrJVTYB/q9D1EdHezghK859tJeIYOf/mN5XK9jpKx1zGxoDk
MHACz7ZJ6Aff2dNhkYP4uV+dfC4BjYFA38J7Vw+MilI3Sk+W5+mEkzWNrpUznxAgckBr9VJ2b5Cu
Z80OP9kIwXbOreO4oYOuWoAQY3P1+eNv0zCvueTaHUCU8b0SXW8v5igehdfjSX91jpzMLwCyODEC
/qUBSfZzmVQIaCsEwaDUOOdf7IbckMostMyYAFGXqM2lMhqbaLHrSfc8HMPkgV0cpB0a/rNYLRxv
+ruBHVJ1t4xZJEXmiaJTUahpd1JlYVrn/pFWwQkgychpNIKVfsDJw9jcVoDQF1tiYJ8gnhu+rwPC
D50vLLlfcZ0aLBAZ9gyPrmmRXhL0aJ+39iIsFpJLKWp7SS5288TzPvd14CmPJ7cyyuLjIdb1KCDO
MfO6tU3nhlQ01kc44l9nvaNN5fqkCM0kvEsWIuGfCQyNRl/hjo/BRn4K7b/4EYN6vVSmVumA5gbz
426gMO8Y5MOXiidoQQXa+zIqBuPZavdHaRb+wBfyJAjqUsg2d4cVZMQYTybNVR+rMPIw7lFxbBFV
aaqbIAHfNPG2SscRrCpmM2Dn0WynkbSkOhyrIBfEB2mqbHWb0Fy+nUql6RiHxwFVUQIHvWvtAcIu
l7caY2BksUEdUe7LdajdpIYcv/wKyjLtiC3+2souFVxUyRFzahbibmw1qA4ExvC2t9EtNEDmwxKK
XEmEqIaYgepHVIdgoQhwNu4+BQV2fDjJGcJ6mODyut6vOjUZFpF96jqBHJnlKxntDCtySXj6XVc9
EAQTcs/vo7FK1mHUQ53V0h1GkYqkMhilMSHsQjkBHSjbunBBtHHQFUChOXUjWgjh/ftPFYJzOpy5
ixwvx7slKPR/lUu0oeuDKnYK/B70ixXnnpzQ2QUWKdvzZ3988tvzB2ykGpJlwL4npGQsbmbcEhRg
TO1ps4lek8OZT84JJjYjq/5k12Gl+bo2oGrQE+zWEgS9EdvjgB0sEuGnTevDXCTNoM3ocv1tQ50X
h65QAf/LrP4X6FRkKGL0DsvW0ZuuDVWrdMRf2XG50u5vKU9EG2hAidCJzGMgbmkci6ACopp1yztb
p+XN9AlOgifWbiRgsOXJnIq6lmAb1VK4TQ+n9kasdOCV8Y5Yl5bISzZfv0m56yptphEP8cF3+UE2
tx82xciZqqAt6/CtGKdFr1NezsE/64QDxbDAH7SBP78AECGEGlt1I3eSoBk04aFivhdrH0DLOIg7
Ie11BTm431D0uFT4za64pHX9ToSD/3NQZIBdK06eoIdd3/7RtRPfkMC01RncznFDEi8VcAhQCzeK
e617BH++WUQo0kVl6nYlEDOjG3eWd7iUCoGR/Yl7cZAc6BkOIFaRxtvM2EcCAx/rXHNW97JaqFJj
lMzytUHQkx3kOeC8aEj7R16BluryVVkUVVXr1oT08zVYa53PJeW3lI4RjgD8BoSGtnqSFoNjqAbm
GnQPtHOYRUx5MFrBP/VsIKnsSppaZQJMhP5JYUwmIgWh13ZZCjPUBuxtmMq06/v2BqhC/0WQWNh6
4363ldR0IjY2YOFaYsxp9s1BgvFTn1yh5D7QOIFNblXsCOvtTJOfjzwCaLNf1/lJl59WzDXomteq
K2H8oPJsaV5qqV7C2YH7xkF7Lo+cyEb3roIZTV5y1qdn72uPqiAJw9E14YgbyfEbWPrv2TEIQP2o
OSEiA8hcJXDD/CO+5uK5tNdaek8LEM2PGVxcH58O+1RyoWu4YDIQPNPMDZcFYu1t3kT1nTqCOeoM
I9ZsLcY3N2EfsX3yuGZvhIiWPktdqh5e36ENElMTCJ3gOz+jlnv3kio3k4LkEzloUdvbhh6hNAKa
Vp5fI9qSYBiTbam8WnHwYqYU73rL6RjuPpCll1MfPt6QtnV4fNUx8W2G4qHnRpoW6tgOygwYlT3r
DdGT9WlA4oK7iko4AKuAlfG/lAALLy380coDdTsDXINtuNAXL4mn8FnaRpqWgNRX4V7gaMRKexZY
PxYEU5zpRJ+VtLHlP3w5DuWeLUsVpez0k/aYhBeMcILFsnPYJgTU2dZnr9/aLUy4JOL8agYH/17X
8iRMyrvq8pS53HdI1XeBxFIqgTMo5r5rZz/ZbaNlI8I+RxFTUgDVcljmVX7wZD7t+da51sTNfyir
lblAelQvEiYanQkcigNuNtjBFotbQokFp6fX5ZfVWxanuLiAvQ9nh0WZOP0dAf1LsV5gb8G3u2Vs
dxn8TkOEMohN65g26WLe8IqclSpMR5ckrgVG7QgWEaBDZLJXY7k4wzwo7R+Uys4wU8KgPnoDLIA2
DNBYE1iiUTYcfLNnbKAVpWOrRaFrwgFJOtew7sff5kvdTZK70jNnIBxlunJU0QGDBq4N04jFQ2W7
cIi2nzRpC6ZKMP6SUzMgdKECiJv0r3ffkwyhnniI+Rk3Xf7PWbA/AfpS8Ce98bU/CHeJLv4xXi4z
fvKBptcv+A6EHYolD4xTE8IOoem5U4H6K4Ox3yZLefIxlcIfRC4CTeN/tMr0p/My313IEUIdBtE2
PytwM0r/Kk3tJ8Bzf5eiVyUNW5+mOAFnJU30c3q1ZwL9Jy8lZqykNc/ZlzbeHgFP/ZyKNCGE4kO3
Y9xBm5EQJhGM+yxD4ac3Ma//wrpiBMCX+qTM373v6WlDVaWOFEzYY6Um56C+iz1su/ggJ0KjKtXR
H5JnWB/OoDIE1AZRcmtbpBbMIoDvuA/LGfhIi6HyFWVQnnGg+1hpG+UZYfxO22YtY3g087bwmkrd
pBNpLY2PwoqQdCG2x2WsCqpBdxoIHKTOXSD5IhRzsgY8B3TM0bnzS+P8aBiJuz7qxxS4+zR0vhtJ
fhVQ79/c3o6+otks7YuQpA2qMdEtMNlsFnGnOlYimuB4PtZuDbSj6yWmo4j0oYF5hb8laOjxtF65
KqsaetyY0qaQ4gSYbOZWejkiUZ9/gQmjpxBbCNL4ifzeUOkoDDTAT+yRWt8aQXX9OIGAkSRVmfPu
drHfk4Dp3wj2its3MYrH6PAXGArpM8D8WhZkXoe/Yp84bK27+NS99pGuaCGOXIFHfqonUGcP4nGU
I6KLjtWTwvdCCDhgWs1JuMm/7FF5bXMwoShr4it2YlR+T3WWeB+q5zMko68nBzjPhQCkYMaSEmPH
p0+geIyY5BGrmd4Gia8ijZjZDSRfYM0juMUSYGlVUcVJohyOwzcp8kq/0o60DXCgF0dy9loQ1zjE
XUYa48qSBeZjWB8/jCTgstVEnyWjoW0qLCWHmu/d+6NGKYNN5BBwZDlwuPx6mHkFfCPcc1VCLSDH
B2iYGGlIWDWHg6uLgNlyv2Pn4anXIfi4oq7E9FQx9Ny8DoUFKX/afuvuy2EcYdOQZ6V0igQfKRQe
PMSdPPnlY29TewmHApddCaD2ZolPm2kDWBpmAD5g5w20iwbW1j84F9eVarNWLjG/50wrUlM+831z
IY7WB/1F99KOfSVY+9ZVDs8e78Ax2bPMeownDgWV9qt02Ju/Nu3CYnxXxJfZ706rkkEjil0k3S/n
wecTMhk4PuS35bbaW6zXK3WCoswhEpEPbcsq1JRipwWYHevon5J0rYs+F9qwo92qEhoDQleEIapA
3Q22RKWXImXJGkD6y4qsUVn61y8mwwhcaobOtsMagSNHZPNurHrIY35UsEAk7F7DES5gPxrB+eMm
jmAkdd+CBL2cDJSPwrLybjTlwfCLzcQYZN20jergSYUoc4CqYBwixwcs62iSC0sjxNjHLY3OVBgB
1v4ECoGtC/Oo14kQKDE+QwsUmMQeSOmX+2a8107SHQ4YeP+Awb5WrmEE0pPoCowrzkpJNLRDvM0B
2Zim+yiLgnKmIEUg607oUS8GCaSPb3z5KFLoYtMYTGxiPCLFLjKX+bzfarQ5uFFp15BjdGkeBKyi
OlMQa9vR+772FyzcGYp4CFQBooevbKKwgJ5C9WKDW3KaET5EjfDFgkQJa5pukuQPJcJfS/djF7Y/
nEjAb7ps0Wm7B16TQvUdwXl/96wSTLrzRvYi7UhIu2oU+pvmCHi268A4Wfk/saDXzZbwW6Zj42uO
TjKkgSAEFyIEcm7kPyswqpVjp8J3LVnqn4mZCkCAaJgoZ6zzTN6nQtM95E/dF/6jtIj7df6SFwss
Pk3KultGumbrfO8+kj+qXgjInYiNqcmplFzx2Lpb8Gp8aN+8JA40nqOdWWzfHqIF+HJSCiHrhk2l
KSCWZOF2Truf8/ZKWGiXqRYyFjjE1hLJDexFnV5uOXhOBl2wZcMRVgBL73t0HrvRDewc3pehjdhB
wQ5XzOt4rIDun4imx/jEJjDCNfNPNYNcghaodouQNFjGsYKzZ02Pbw+U/ZrKuE36wOwapz2qMPcR
mlR54D1l/PUoxX8n0pwUOJTiLy5EzmrOr+XGunlr0V4DCRQBri+xAgnwvLOjZmjWdgqjV95V2Qbi
yUDWSh7pZi34Km9outWX+ewa6iH/a7qawfvcyciB3pFaHOifooRlsZ4i8eLv0DXJ0eVfchr0mxCz
AvY9sUtG8cGr9mj+DfOgZKT90ggvQ4bLvWx/lxbBnCv1nZNFhzzn2teS01xsFgzcVxC832TPoZDk
DkwIDfGH93QaZba7zX4Yx4efAfW/BfME3UPbo54g0GtInaSUNm0ZyA5wPlqNwSx/YmiOARHzcl74
+7Mqbn4C4t7GfpNVrNJG5kvxvZxldCTkchUXMqEo+Os0WYEGBXhpQ3yAVUeAwzZRN7TbkPVaG3Wn
sM/P0430KI/3yKktco3PF5I0M0FIjc9CtMHAXhMGBczVp07RURC+fwmeRpAKk7byFSdiKYpJTEbo
2Dj9ze6hLBfey5DpuL9FBXYMWLE0C69jFdAGCKCE0Pe4hD5m6zcO8ZGk5GgewzNAoN9JMOFm3eoY
hRsVbtA9x3p/sMaHTjFhb5W4uRAwrGX0Zkj5CkmLv9pA/HDRmjzo3p3gJv7KSkqtAj9v7xhig1XH
fmsj+qYmxMWTpmjRBINk1y/tA3bbvwf4oJ5Yb0yyMy/p48kCPcRQF7hq83wF07b8yVCfZCw1O6e9
TyEdnch3g0yjiq/WN9AlbLR05BIFGl/Wc0/PwgRFLwP+vlueefRtrv/xE6Pbeqv5G1RzKCh9NLO7
A3StHr61u0q55KHNbAZMcom0zywV3EVwzZ21kwVikQFzJriFDknvj50212gNd0ej8XDAijlOSGsP
8+YLxggf37WL6OgwHUxNPmH7sgIjDBkEN0caG2+pfMQmC9n4vLpNfPpyBZSykoOwn/LdlDFLR9K2
V8XgtRyco3UeqriNTOfSKtliPISIsnNMyuoPZejGBvPD8Hc0ThfTvppmYhZoDSRaQrxy37XcJAWC
S1MEF31an2pWjPvEXp2WEneFT+CX42gGj6adZAP5Y86kj6YQbUGoph7M0Vpyc847EhInS9fTLsDW
I5YRnKFt+pfaZLsphraSzzso3xyiyRxvAsxFrLXB37kGTMa7vNmUMHBdIDOHrkFZeloTtbmzomM9
L5BIJgewUe9yI1IzS0NrMtdez6s72ZJKGmus/piNavG1jI/jQM2TShtOwxgmHjJfsEEX8TUdcUN9
VZP60d+TsnTRrkXLHx/uLU80EWVaCxQ365T74YDGQ7ZhsZc85YBd63aKymYot5YH4k8HTHRG6p+/
Lffafc4G16GEciLBJ2amsojqUfOhI2W+5kc0ZqxQFtaIwC4Sb/gEc5f9KnoyVteWO9QG0pBuBezh
hub7PXpU55C5ruWCyizg5FHLOlXqaekvt+CMWBhYI+/i+BclU32+wJyWEKpOc7YuqM9EGYiRBKBh
01KaldW1H4VycSD2V4rN5bgQtQooU0nTmLO1sDFtXFq56h/VgkRjcTiwSA+d/bTqlsY+XNw4HTUe
gm0nQgS6zaLqWPB2BUKlqubX6HV0RudIe1gcJcHARkYlvVK8UPWZcwLpl5yROJhP7mdfdu7wC0Lp
rvkecmMQnarWSllsHIwl2JDlCFuXkG/Yo8ahb2wqI5ek51AHSX212PTESkoRPGAg3VGIggpCQcFd
WbjTQmVD6oG0vcoK8pd3Luhs4Zg9Z7V5bgg1jILfkFPoXOi7OQk1VGPTgIi7CUnXihSWus9cuiuS
rkjCBrpcJFPVwhZEWnSEMsa/1x7PBqEx2QB6bt9u1cLy9mZ2yozCzpukdO8wJ4WMM75znJ11ypno
Bv5O3qZ5pqHlZxGpZvs7DR6KCmiPYW8keDekZxckf8otULEJAciaXThJC0wuTOolGxeKWTAZqqiB
QMCXuvlRA7Zn4pWCMK2XKkgirscmjm9mye0J77pmfG0c3jKYH/pZM/QgEBOQozsLu2OXIh7LGobT
t3Ar9yKxKGAoHQoBZVeknuvb6m6zkxPinbm8MxzxVf0vRpS1gVUc/xcU/QlAp8uZR46TEbpOQNg0
BIqZsfcz6DUxqeZhi2MhlDZmB6nfHlS6HSPUBLO0MSLrCln35ov6eCA/kQZS/ZiSrsy9mfm5lmCx
NfSgs9D/0qWxkIGpHpSBLEd6RVTYzpOLpZviwRmbWit1BEF5F7VU1LAZ/W05yovu7uIXRUJRg3iZ
ze7A+jo4t9cHK4Necu725Rz7r5DqYBcNYC0+CDq4ZsM2q2FYjVcCwrCmo32ROAbB7xRvcbUzUKkk
jZd2uyvcL4Ah9mQhpiYbg0sAWO+QfnE3LFliCfFZXo0RxcwCUphAddj/spHkA9SDfGZwHAO8Da3S
d6kyPniGvQ7rYxkACA3XC9HZ6mYVSCQmm7BkzULO3T2tA4zd9viR4KzFKMtzw6x+1mJ4DihseT4R
yYZOpV8IcTSKI8LTPwvxNjQy35DHFEUepEmv1TCzxjxRoq74ssttdByXj60AUOxPr/F5lsZZ/O1F
wCdPLjZXbwjnq8lvWRBkX69tWco+PhsQBArGzktyqGnDf32Ba+9MKmmvtRPdA7CCV2+DhKAlAW3A
IgdTaxhqg8mPpT8cXQcedDdnnZJA7y6o7HRjwDAVB0ZQMuc4KGWMtol3uwJJWBRtEzMSUCL4jFC6
B0m4acJbWTignXCbwJalQeQZjnqKdOhZ4wmOJkuYBEFrLvNdkRAENC1DCAKUXeYpV99XIu/qELQg
6nT3U2akDjHDYCI1+cnA799AtSVqmjO8A+Ewx/R0Sr9bLiaImAWpVzzwA9cvHp6L/fOscVYNz0QP
7nI9XbOhHZm69b9QdxNHNW7qgH6XNp7cfMffpbCuLZthYX3pCD99TGmdzBRX1aGY0nQHaXgGiFHv
ikA+Q4NPD2/FxeNRV0wORGRohqq+uJkoslereNLelW45ueI4lBtYyWFrgbgpDVPl/xYJdiK0s923
KOA7nPkuOYmPhAHkWMn9P4desfZtpOmk2r3J5vZcq2tQQcaS8YIReJEKXXfHf1GsBpDR6MVGors8
F1g7/VKbtGgnDYKxHX2hekaAnodjl6ubNgcLK/w9QMbykETfJmIpM6IHD3yapQhDGAAPYxMu/ZRv
b4YlWZB2+ZppSaN4/gEFmHcsFZWUN0ANJY68TwMxUhzlQncxFhRmsRLnLNXFJnYWurHKSHwrcdwz
QavJOMFrKzEKKS1nkgZBlNCz9cZG6fcNnklqK6xqIh4+GTNYp/sJStWuCwd2yhUjhjHrxz+409Ti
SuPksSKr/93Nz8vuDV/WUiO/OyHVmBeYZWpuSr6PUbSgc5LMjipA7Frxc2GuojnrAKQxQZ8c0SOy
OX/ZhUDJmOFCc+K1u7WVqZ6KsT5KomsJAWUpCJ5DjPBp6GHhGAl9YCt0XUet059w/aO3PBBNpa9l
amBFYtRrTH5GTPbAXwgmzqmFkffF/BE3KzfxClyL5XroGD2RfViaNJsthk1L1TljtcH6jTFZa/wq
Y/jtVUmBYdNtQBDXT74wvV+gBXe0FnNf1DvwecjXsbhFbAGA8YS6gUfexRYhXK8tCmXU+YL9hRo4
lOqVnhpLOIg8uGhcR0XLRulsuj8fnjbTuVI/balkbgiDcO4mih06WDnl6NJPB+UTFaxydtChkp+b
sYP1yq5h9kVmZox+3tljm1/OnYjbX7KPXkpLH9ELuz9V6lgfV0FAxL4TGPWJyQcNh+6fMgQJc4MB
m8px8smFKej6TZVsW5DmLWuIy05fH5ZJVw6AsSjhuHkDTLt/igqaXgwX5+FXVyQ0L40WGqTCV33K
Osdx8+lFU1k89b0LM75SWoIgyzGmDCCLM7xoZ+GKj+hb5pKtfBjKKF4bWpqizU6XwUINDwKKKTb6
Y9Odsxac8LKShF4pXbLvF7wfzYAueT7xnE+RQovo40elPAVQ45EwnOi6Dhka5hgF9+UnmdK/s5xA
jVhAImVNSKLKUI8s2dD0wQNqLzGEf6fCkJ7Ccs7D+bTwRU21AS09GbTYqk39z5so0+Xn6q+qWfh7
AhJKUTF0RLeDMHa65wTTCTcDijHyQAwQaiiKWXKC6zbHf6DNk82+E/G4iBlr6p5eLI3Sjv1sG6lI
M53gU4RwjlxMpCMi8QXS4kqpfb2nKv46SapU9keAYhYDLNX/WsHblAIoEkTg1Kzv+cf89Za2Lf6H
qt0YPTvDuKzcf7F35Yy7YD1czroHVkh92B44ZJutXAfTMDFdI7Qae4AtdRETJcM/gq0uQ6M2hqtg
OWmnMiH17U3Cu2Hbs3Wl7vIA8CjdpqYi7iEiLLOkfxqEO7pjQ0rRjYwqgLBFpWn4LDb05NDKIAD/
fc8OtWcHlFhgOlf4QCkRQicFiXZSJv8kqx/lM8/b83zbfdj69vPYeGVpxo2zwAKhMZonoX5WfdQv
ChOTXYr0OsDWV/MREc5RzrMzMUq5ORC+N5PVHF9lU3JAYFcKYdxHf1wjLL9sp+fhwa426qogy9Xp
eeidoJWvx3RyzD++OplsUxy9je3r35gc9HpdfbOFByw9gHDm6A4SfS2jDHOFxNA43rLlgQpMpkq/
3ANWCgXccgTPR35Cn6Al4In99Rh6pFE/ifL4cZf+ftOQkTd/t2qdGYcMmKBeruWZEg1hMtwCXUe0
KacLxFNYX/QEikzhBJrftz7erBxsHWMmU8vsEynuZV6ehQ85hf8exszXsXoIq2lSkmSVZRP1E/Of
nUb4qQbaHJ816vr7LWr73GB+RgGH9jRDhKEfdO8bGOefOb9+tA8S86ycTgOzFr9+F1UighvnI96P
OfifgtSiz2Y/naamk/npWd3edt4MYg9R94Ripd9fHmHzS7eylWxSVjcpQZHVcm0lZGHnsecyr44r
QZkmRy/prbuQAVvdmpUxPBmKHikw+HfFSi6V/JWJeHoiDARyzf7CafbW/pY22Ec6Xn445ceRaYe9
UFwz0NoYWbG8d7CydyWeHDaTvU/nIoBivDCBDgRmXravn26aqY+0o0hZurO08e5/8/n4xnARoQ9u
BJGDK3piG0mSRIuq4muaJUwXj2NzEnYfbXXBdVqbVBRgZhp6cQmi9MJXa1X+yUrHJdaBCbt2++ak
Bz4e1N6Mc/POfb9UrgXATCV4UTnWoPeU79UVqby9qMtnpUsO/n2eoTdiYYB8mKf7YcSGFp3oOfCC
vdWXT/UcVTbXyOMUdhAkquV/Jt5Gs1cTlQyXIj9SAEk9aw/6IQBEM4lAst77ms1619rfSHEeiP8h
yqXWUnNrzRvX41yj4SyYqwR63MJG9NlHs9iXTnlmtPviCCFsdfVT4XA0acgvtSprCM/oNfniaBZh
8L6lTCpD+In+kFMRqQCXH1f7vgyO/JYaDoA24InO5pas2eYmrvMhQMRC4Us2GBMUc9NpZQwVjlBp
d9aotb104MMbgHgBb8C+EMQmGD5ilbHVRuLZK6Un68CLlXZfgqkLoiuqFsDHsD+i/B9FoA8sgaOi
2UM23BzCtpAnWtYVPMwqDeCP4Vxtdb596GpYnzM+t4ltK9KYJYDzdhbng9f0rZNKtCl1przUtgmz
uDenE9tdMQjpzoW//2yqMugDQrdm88LHqrEHMGUAtP4KxFHhUwRpRD5J8AIoWCEAJ/rFn/x6HzHc
rhi9QtD1exZes62oCireoN466IP3H+sNxgyYPDy4/KI8FgXVkJbU+KujjB2B76cNAnfjRQ5CMJdd
nhbSfVcrJKXJCwSr2YGD4ktwUJEzxCT+9rSZkDFbJKYdqIAdRZiLKvnVe8xw9UTQ/HLq0wxwsWqM
n+1glRs4cwTDifxCULVzxp0PUFepW7lxyr3xlAuZ4wRRC3Rf8a4JKXXfsJN9bUu8Mw1VH2ZjupwV
h34fmt8xkvlJmIUuzzrEW+QTsLZxE6Gar5u371d+9n0lg0AJqIYH3LGk7HMB3GeorN1JS5edysHk
cXUJ9gzca6gHwoCPmnTD64F5xgu//fmACu+NGP7FIlh0//DSHcpUgfw83eFHpdviRcZYojKAAZmg
JRf168jQ049X6/VERBT/7BfnUuXYEb5ECEKEHA9G04D4vY920SpXT5BR7Z4wuAgHwdhDNaIdx/sp
I1D6X2rhWMY1QwTq8XkWwxcssxTSqZNoENk/MVhgZOzlgWsY7K8sVzd+md4Q9KkmS/tlIK6nF19h
cgVREy8EgwjD5+F5c3chUAZUX7jgUkJqK67yZO3V+RXCk7WnKqfh5ZEGpz4+gyn/fzbiBJE1X+x+
d9fJAU5LBv7rlxCYG6d8DlTpTPdV3X5SdC1z3ICfmOrSkrU0H+q7t+CigH+hIuB21DYjrLM783Wu
9CeQGdKSuzbOlFaXZMuYr5ZXWFrMnIkihP6tG2IDVFpPFghKWuKTvBxirtLarQf/QE4euuwVDMkt
Oa9mA98jZv9R4h6RrnlEry00a7IB3tmp/3+rE6iUPTLR9XjAbgR9+96ZvHHVmDFnVfTkSQWTGqTR
VRG6/45Dtn0tvYamFt5VCW7dVQuyDZiFxKHNrUO/Q8W3UC7Pr7so+BvBwL4Js1a6c/LZ6LeuKhH/
RXvvmksSqvq1HBTP18SALumRlQAir9kw48h2ENZtltDR3Z8Rg0mZvoJ32e5USLDAvY7dmNW24exV
BnUlYpxZv+T6/+ogGvBpl+Ld7wRr5jIann5kTDwJai5dZC1d+agFf4fW8AWyCHNGg0bTnrPHrmPs
15oV3yudgrD6F8beqIb5+20W1xHCo2QDEuG2+hH4oH04WdxuWzs6YIGQde6b5vGpDPiKz0qpn6Fi
VsnUMneJ32IlGOfxO26gV1jA34i4YoNmUhnxvXFeYHVoKvMjsfZlqS+9RigqNjoeLwCynITcPLbM
Ow+2FxcYPLQBqITYcJHL92oW5DcF1bsjVdYOR2v7XMsVwGwKrF0uJk/SyvbU1xzcyDwnN1zxW4WZ
SpP8vv78e31e/EtmuLZkHaElpvTdtyg2ut9UsE6zsUXxp6yQkLwy+IMqdZ8oOvBV1D2bAMfY8g9u
zHgUD9BvaOqKwuLhunDs55G6F/wzv5kgs3JLouUyeGCPM1bHtbsPb9q7Mq8JTvI1vO77xYXog53K
P4sw+wWm6tXni6/ToQEDXf7pYLRZMYNbrkNm4lWzBUWUc49sVTSWG34KmgJ0gxAm6fJd6RWVgJ5u
vyxJuHt+tN6dfXx4n2kjUIwedY59zwiOnpzGm1WGagffUYekw6Lneqxcf5vsZEU+Zn1CvJ/OEC53
NILfl2DRUU6Fjbqx7Or5bJQa0Hasp75wjaxTuqA5hGrq37UR9l7tcYaRidr5nQYsZpTXNB6tCLsG
1IJkOiI2Fj/t25t9M9bP0eE0SdG6WOWzo7sXrbvw+wtQtkorJAcq6+1HIgKERJ6QSCcFuwPoOns5
j1qpAlWzNdN426PesA8xpi6iHinILMSRnsF7mNGhS7aqpsBypUipAhMrkr+9ZL5tK525YGxPYoId
dSsEM53ibw+LjD+oPSbTIFPoPEp8QD8t3BfIO6yNITpVhCj+VAqxzC32+05vv89aJGDmylxeMYad
O7Hz4EX2x+lzpqCRzExumJDGWdpGj1bROvFugf9Fksc16kHzqy04pN1pPoMYByo7iejeeN0Z8PeJ
LcG2RBoIEnYwfVS5M1BldL4M3CHnXtjVqifHFADVOOUyleGg/YlaeStfnVxSc8j5IFXSgCbcyLjy
PbtM8KgSvr21QqR0pxQ67UEZsddeY8fVlGjXX82svGc7cV0iHlN0mP1k3hX4+4ZEwEskfelH82J/
GJYH3crCmB+1zVSGWAA35dRJL1GU1RDhUcxQAQ7OxrzR7LRGuBPUuxOZmyOesfZDTImpwNMj0/y2
X4eidnXBLbzZjQBTxBgUD2AaXkHi2LHEPUwHVM4CiJRfn73s8XOTpTAu8w7fLELo4cQ6BRv1wKUk
3pvEMiJII1WvcTVSe/WcWpM+NX10ZeCcUDGG/6sbRONM/3uofB53eQV+nQn86K55l4NuKbW7Orqa
vF5MXTdduwZ3kWgb7/8+r3ryXa4QYmwJkMjHw7jpBDZTIYk/1mzD0NMadXNMjdUeVLaszxc3V57G
ExB1mSwylNgDH8EhIKDd5QB/vaU98SvOTD4BB1iM3KAqUpNPvbfzappWuLoJcrnbGRUorvAf64HV
hS37Lsj6w4gw8TLebvCaLjSAYs4o6puKwYMavfnG/ljnpJyon/zcpTOTvclgWmfSTC6ta4/H76fb
fW44EqVg2ol31UDp4noNJ/moDoFyf+iP/Ld/gTBAAxQda4uQ4jvum22iOE+jdhjCrbqUCvrD4IkW
jFUxeYHLdMbbwg/Sa3ustgu2UVrRPpNNiTuoV5jSkb8MRw+mSYELEU+w6JO5P2xf5MoCtLjPgOVh
+vPXHGCwKIelzVaopEEKylfFaHqGklhgLFuTVl/wKvxAh8ketROVi7Q5hNTfzVn0AEQOKD8MbkIG
Mu68KvFWOKGa5/HX/t/K41EYTJauelpwu0FEzciEYN2p93XRDe8JPmGHovHRhWs338wT9k+UBpK6
bceqE8q0g973a4ZMJA3b999NnTzBKP3PvEUXZw0b5GCMMsQG/OGlYM38oluivAzsxXHsVnRGbfQa
1EfdQBHHviCU0cZGC5/1AgFoMghjPhwI0oQt1V0u1V2kop+P6IyjCp2evzSELthIJKnpOaEZMxgQ
1UFfFEPb+JH0RKcX8EEM6FeUHEPDvtDtvt65xtuNNF8wcSiPnpcEV75zQc7thWMPgNccfiViNHqC
my15O/NW32ciKzBNYqbTWvAYjx6JFHpsmtv3VgV6btZgQlU4qIHPAzjf+sy1eZqt5ZHdOvoPfBR2
109+CzqsOtAVA4bgXnv1mDFYCakAp6v/VeUwSLMUI8wxd5JUeR09mDfbyXNZMEDWnHgPINIoG49c
lgtxkOQTnBhk1zuOoCQajL9bqd6WZRzJFArBQalQGR6q+k2DB+d95w3xs8LbX0DeXR+8LMKk1Joy
Q8N99mxGYVSM9U/zJ6nTYfdQH7eavPcrWH8PGXssTS0fSyMbOSMZc5Ze7shFmmxRcEnD+j1KTV0X
A/0p3R6lt4XRwRxJuMDjlM/gDto8xJUAR4TBOaGW4jXPxyYMBEEe7N6CFqd3nMEZY/X62du7lWCi
2FIj5IDGVL8FURMs5xEtrOLGXULwnMOIv1BMk2fDaUUElWI3MGWeXWZbrnnCyYjTOIwWJlt2t5JN
kOMhWlBBA7iQHRecxsS6CuIbVfy4zT6+I3xewde6Un5WAdKwva6jdwDHsfTD1htpgxJdbHsx+FDM
Gf5JO06AQq8XYQ4tX9OuCA+0f9kN1Q2H4L6LcDzv1+i9xiaItKayzMUfMaI7vN5TJvplKnOcVrWR
Y7z7Nh7eIhHFyl0vElAzHjHj/bv9Hr6c/mWbi8oBX5FYe4ZFX4dtmKUCzbsyH2l5jOTzDzF4DxbS
GTqhRjXE/f8MIs3zOB0sNn6twKgwIjsVZ2LL0w93aI05O37/h9qYqC6nnStfjPr/k/im/3u01eTi
kAKAz202dcjse2HJPzoAHYD88ldy6axzumN5eCroVOG2cRT/kJlKf7Y/6oKOt1WLtkOumWdT8gRY
+TePI959iAf4MiUKzcuZbWG4C+V2CN7pkrFt3c1DqwlCGD+td7uVxJrBN3QO5izH3RvWiiTkAqkF
9NIujfCJYXeXvd9HvHTqWiESSMOc+4M7B1dGGFdlMIWKD0lq6Dd82q+9Q2BngClJ0Dewc3yybV28
BkZdGbfctBQQPtAJ5v9hURlmgaD+A0bo24svyRxyYFKjHe5j3RWylGOOIavwQ7fcQJcxPACbxXDd
ZzA5FImujMvhFWZ/z05RvssyWNDnW7+AAaQ570ssLUjKNCkgoxDg769sPuebz9EBh2VL2RQklk3q
POar5+kSPv2LFwjlNLN8JqqlV+rQ7HnPgOr5/XNwrECGBVE/GZZjwN7o8NfIC7Ya5Iy5vkkB91f0
F3uy/TbZMMcciOx+rPNheuor8O88ShQbCPuCWKI55RXZnAz6g5TjZbjX0mPROrLZrJBVO/PC00JG
uebYrWSRlHYjHHFozirssLw1ASnNgjAqPltX1EoIQivj295Vqc1g91qYwMM/tR/pW2pfkbuNeeY9
Rx370kEBNsBeEzTSbRc9GT3+0HG6ouf+f1nhI/WEs2y7w9wI83tN9KXY0RVb8UVTWvfhth+DSWnH
fZV29n/ctXl5b6wxVYQ2QcZ+CpCjPeGvhaAe/0UfkhYtRbrav6f2miSNOa68plyQg7T5apjzIlfL
Jg3h0GKq3AKKo0ixhiy4sTDPrDfmfC05jNniJrCoEKYOvexXnFj/OkauDfcD5d3eyVDnC5gZNuG7
zMy5FrMqviRlpC3x/jXSufeBbf4ckvq1Sl6fJCR411ZyVwsAIke+6Ezhr8mLdiOqJHvS4X8BQZcT
eXpXoY9xqpuID/gNUwAzMS3CgjXuC/KA3bIw6FM3lJ3Hs1lEtS+9Oxkj50uik5DUCIdxUp2NYesb
J9vl7uB1++qyx6/JKpzSUR6FaenrD1qvumMsEZqkYLnn44tVek2rqsn484m5pqp0RVI1rxw3YXgZ
DYP4L+qXACEsGEP2gM60MzFTTY205THns6IzBA9TqFkJkOQ6N+n5yTc8YvQfT7+WbVRW0HU6p1Nw
KtYSGI89RAGoFS9MYu/xHCFfr2fkpamlNcBgULXLYP1c6LE1Ww7WxQ/kEuF6DcZqX3RkgcHM7WBy
UoFR57twk1dnaDDwpYSnR0eRjo9Ttpe7hDoeFHdu2R1sJQGqHZU8Lur8xSPCFLf3dxbt5QHZE8GD
k8CXBWlIs4BEfd2j3WAXuVJkqOCt94dYLxJwMdMtGxnQ5BYXJUUbBVDKk9/OXPrv4BM5bqmBvVUv
QQE+SKKxCARVHfqvCo5E6N2+oGpbNJwH+zzC0mHha0W3GDMaR+raV0OxuG5AoP+ZaUMGB155vpr/
+c6WB1ZSy/3Ac9h7QM+Jgaf6fvUmUZorgErRt1gdKsNpOSe9U/tZwC74n9M2EQM0yaGuRKlOP2h6
rMAt/3rdZxgnhm+LthrpOIiCeAceJ7CZX8mlIRj+MjyfHiwviIT1zmc5RZzYoRNmSTAsbiVreAkG
NABlHzyFfluaf8xtBux7eAM+PW9QMHfISXBIIVMMht68nQtNreSp29ba2fEGVmu2A8+ckeOWvVEl
Ia5GbrA73jGSwN29RmDllf5Vw3N4eKPI9GPOLOVODWhsaXOzehUnDShBp8tZIBEUXm6JYF5i9a1D
cHqAcNJgpJPFczO2TnFZOw4pzeXe1IIgwIpzWYJ3rpkIuM6A2CM2R4uQBO8aoDoBICkxlzYAUaMp
e0F0yXm8zNgsj97lerTU4SNOBfE1Ha92hhYyLMPvDv+jO2pqobLgY520GcHAoA17buuHi2WSlBWK
8dn+B2+XSf4mVrCRRZ3ukKZB5BvCFuuPsAb/oYWmzYdzIxT/zAtMDa7T2EWoEkOl8MqePFL73UN6
rCePgbQyPbgJ9sXhHNTubmM/fDsIk8QFuIGlN3BiiLsSBVB6U2xEW/N8xg1tMrVmqlZIkA3sgeos
t6nV7jY/rTNFhq7afexD+zbRsnMmSLNYsgkPRbahK1r+jo3wIHkmzLjVnx9ykr7Hfb7GwR7PDkVq
WPiBUSBG4eHrM6yPXLocN/LjxfuukDQdaROJK6+W6BHLbYbnNmM34WI+rS8UQKqRziMoIhByN1lz
YqkLaK/GAljmZVA0q8pDm+/m6B+88irvbcpoglgPZf7mgJ9zFCUkX5h3fZbSJg1vNEK7j3JEXALf
ExuCxHUPRF3fSEKGPAwcHdwt2CrMt8tybs653mARJbRgcOZj8Ii2PvhOU0qxSR99DVoV0v5boDp/
Z866PUlhcbfu+jQ0Cbu7t/doKsyJKOA2N4aM+gtyP6M11mh3f4nOz3QR/iFzkGM4gH1tdp5FXi/g
NcoSjIMmx+7W93K+aJGRj2gpXikWpbZDZlmikNbMZ3KHwxDwUsdd2aC8DDSXG5Xd1Vpr7n+03K66
Njxu1qmVwA+LQQeXLD6li+k2aSjCuI9fZz8tZ5qCPjV/OanA50/JpoLJ9kKkaZaIwFC6KkzxNF1w
lxNIjOrEpa6BNkI+gP3G2mDHI0c9HcKtypflUf5/jTJOxly2NhzdkesrniApBFLeUX+OIuRdlf/L
NT8OOf7CNoJDkSmIUAngT0kav247XYKLyEuaM3WC3JRnUq7bZcUvtFrK1zVp2BUnnP7aPmWH9y+T
AFXCoK6EXpzbfVo7xeNCqDTrK6FZ5bzQPJp951Od49/6EDJr9qg4+mq4SQ8+Jy96AGUcB74JG003
IbsQ9c1ouz3BAvXXzj8LZMDbk1s63xtCAPYlLESxp+ivYno0nuLWjDcsBrWiLez3OXDgfRm2KQIc
gE7b1Ab3ozcjqwPaxK4/2QCpWpzo31fUSOZckdF40Mf5jAk9Dr2CqX89AyWgSbBIvQdZStOZiN3Y
otk0Fdv5Jps1xr9Yk97VkKtSFz5aNueYNoSCciXVsxfKGG9KNMBwKFtgaqcngPW2nEAf3N48O9yj
HQsu/LKYrS+wXHQhR3pXWFnXjiESuUwqomr7WRI1W16ccIK3GdB507IM2PtpJ1e+z4lxZWis5fXr
EwN9YmsJrXSbNbshdMNu3lwqzLVITgEtrWM21ESpuss2XHCjILKjoiQDgvkvZxKjR5o4L8un759C
fT2ycDLTXV5dS2C3AUbXARyd3E7utl/v+SU6LetqmlSkYURZhAXfTd/VF04qVqOj+a/T6lEQat9v
3uUAW7mUOnRKdFEX90w7ZdBOIxN12HdIYCF/V4QrqPP+TItuM4mB9Pb38YLweM4y2PdxmIAecDOw
kAZvlQkwIlPk0FlUAWZYSwqh9KtPxygFJERTw1SRDp0uocERCaxOmYhk0DzYE+j4P81neEbtYLIW
gc3NY1MsooDJwMfPOAqIa2WEGoI1W/CdpqxJCUfLeg7q62iHAJ/4b5TsavfTS0cwTw/O6JhCv3fp
fokC1LhEX0WsBw6ERi14mPaMf3nXyshw/AvHHgCVrgg2+9mMavaOxL2rXgKa3i5nXRkkIZKnvvJL
QhkzdB2lnpKr76I6zEkqJS8G/10gNKhWUIV4GkcgK526+lIdRjq0J6NMX2ujLJqDW80GgTNV0E1O
JhDXOCOkCgKgmuxdx1zMF/yxtun5Sb69uBZFNy2o0oB0stP5KZzZKA/9GorZgL9tCrme+Q45E1VC
dGFPSxa7H8p8OKH7DXX1sRbePczL2XnqU12iUj9RIHF0HbZdcMxcsDXwkVpJmVsZoA+buJfvBimO
x+NrTkX+CRMiiPYckC3BtFdzqgjk4hxLunua5rTtmXDmW+e/WOp1VfG6VQe5HFJyjhE5LKkVNrxH
0J0tzmX+Y3NBXW6UTUIvYHipGrNk9s9NZzSm/mmDJQFTUtcslb4oM4TolWT29hkNok+EWBOtmNBs
Dxq+LXuzLl7TjtiVZpgAEG1nlZR8+xOv22m9ZSPVhDTcbQbWPYW0ZNZ66CMJy2VBd4mvHA0J3bZk
vE6j+ugpWRLJHqD0D9gEkrg20E/5+xOT7lXO4elcmVWlPcQeAzS6x+oYD+PIhZvc6LW+IHt2mP2h
9fAAuPbZROsnXA9/aqwsFeMHuJ1jQLS5hmCQ4niBis7vk9aoAdQjDjA47u1dxoALk0vwmWv2cWdc
vT+YXxS45rD+QenaVx55WRyNJGftPoKU3udN7iphqjyUUv6LCYPqA3VUz1V3SKGKdfk/VVhyvla2
w/UOKDosYq5EdTRDQ65SMxYr7yJlytMNOIsqJi+v/T0phxC7Okw6ae25azYotiMlnSaIttm3EOqv
cGaHesjhz+mXXrsPjgyO5Te9LoeifmkavX4U4xboJyv9twDg4sZq+7tHUn+m3iv1Egd27gd6042z
H8/jfLDY8eFTTvwhuQsBDeC6vfiHnfRTk8L03T65X6H3Q400OCiOfWPSvd9x8sCjRl8lhClowmcr
T2RNOp6kU+Nk/jNsEWSzhZMSQPM80GBVj1dxD1jg0ZuYsxUEF9v9ePdoXzi+pOE4+3wezpaV27J0
oCDX1d0BbLEdTz8pBuAO9jtc+T1x+jTmNrRH0f11sZP9VCXcoMOFYF/H+vibNyq4kGHotUO1Ak+0
mu0p7NiK52K3i/7lwcnMLuTZeAOft8hx7crLu4muC+Z4MGNYpWaFqDYiWXyQDpIgnsKNdsY8UV48
m+lIZG40faFk51tGqumbOZ6fm43Q+ZuAxsc6GxM6sivzwQCetSBTbYT1ygWnyTcaH+k92TY8IBJu
N5cU/4DTySqqGYRqDSpjKzXx4uqlsB5eY5U8B8wtFnuefhVs4iPDm6SoIdXRfeJiROcHQFZuEiuc
cx60KLGfOviX9PTWkhws0ocI6t+spAy9Y6VES6DN9e4Gzx+Ao3adyCw2fdDyGhhxrVbtU3Vpd6Gy
6S+Wxg9VulhJTKikRKjjyubRH9w/tsbYaO6MXfNr4Tx9IBPafVJag0yrwoIFtZmgbrBwj1AV9Fcr
vCTvyceWMJgg5RWRxy6CxbWxDy788JfWAlP4+XDt4PSeU/tf80GWjx6oHt+Y6BoLH0GV0ShKJkAG
BLkSzMzzLSPhlwIzrDpPgV/pVj1d6TnRd4az+6uVWm6QLm44dxRdwFGxC9/bQipncVstnft1YRAi
kFLiE8NCygjLv8yrGR0rLhS7yh8V4zt0U2OrxuFr2CdfcN8vRNaz6XwyZ4+62Eh3CwipGJqs57W9
mvoaKr0kMiHHM1VqokDMhUxCCHpRiy2ImEIcgtxQ57csSMZq/G66idWt7BRSVTD5/mCqhvp1kfwf
v4QFwE6PYU3ThluGuEOx4fr2kK87dR87CAituBVcmPsObjft++gSMmjt56NsSQXYzpoUbDE+0J2I
LG8SqDVGJDyuABimGeaxy6zShFXvHtHAgSEwDHLLqxXl+L/b4Kg2GGZLdbl5pnCERBkq4cxqKrjh
NvrjdijJHofyDZ8nX1Jn9sHsnWxDPbM0GC0kVMwH09BOvX94CBw+93bmrio/eWRzrplPjgkWivE2
Vu47AtDXskKUh/5xrhlq+F9Us9tppAyb4stJYB4476yCfPu1DL/AH0S2CIPo6rAzd4chdM0LPx34
7f22H6hIeyMIrFzfwKhtgUsm5fGFHIO2ZqfFVfxRtV5LYzn39ych6pSBQEeKuzE89r8bTOdz6swn
P3sg/Ilfu+i9Wy7jyFbRGzRmOOl/s1FHp0ajUtjeKlIHKYQUSV2n3JbHYC3CjBVkIaw6B7oHFTTr
hx6wK+VgO5JZK3AnGkaTKDEOwRcaO690tBZKfs4MXV3XMJ6ALLa8fJyU4q9A85HieoTV4Z43OKLh
v/IqyXnrb+BicaMxfkxo1sbJkVBQlLqdwaZTRwY4tpBFW6Ib0m8jL7T/cHJxMtZFhXnMYuY7pbC4
atsbKpJtpgCx+lXOmNRiK1q2ujQAkdo3zBpq7UHhVxdQycDrGrGsH8t82ujgVWDZkgxc0mfYhWco
nIRX6y2ukDljq1IvqsJyBUPGVwoTPo204vnp6guF6VL1t7rv1Rcj7LxkFpNA0Gatk4Jfvm48G8EL
X5aqIrReYus8s46ri3rG116x4rPFxdmjf9bYN4jxBqM9SS9suGnyiA+kInAic5YfQ1D+QfPL6Exe
a/gEF/BIdR31gQaZaysSoI48yePnQ1oXceiph7wBPlHUGL49qC3odGqAVQ9sPA4NpBUn6QyK3iky
gKTWomZrtl9zmgGUe/OTlwrkBt0SmS9eqPopwl/eOUjlm2xkchNbOvybsPEjCjZ2/QjKta4imlcC
2ZSqppy0A0fja29NzDAYE+58MLuFMpDdGzki/asBdrcOiFQBCUs0s1AimvzlBORfY7pDajGg2arW
6WWfb9zeMK0X89ACOeivdlufxyKt1/j/Dx5K3k702ByUS+FoLuJlx+GpD8l74DbYJIGe/R8LDpTY
B9uPaP2rdsLvG/lipzrRqQlyuUPy3JrvAvbeOAYfpE4qGHTPkl8U2bS+sgukhJCE/YYFz71Cn8r1
WyWyhw1z76PQraduEfL3Ff2E4isnriQx/griprxtzBdBYqu5JZKvIrKrmzBnRcPtyiV5r+h1qBhR
hGtmuBDgbP1a9nTz04Bq735CCKHpebwv3R85Jw/93fGEcFTJKPeGNK/N638e0QgRcbuKPlpU5pGl
/qer0bv3kiHHyAPk91oCaE8NjLJv2/i4qKLrk/7nFxEHzQKyfTasLzinikouZzZ7XHipF1FISyOJ
gkZtzHFMoivS97pS2VIwu6oNWg15MRTq+z+LHycJoLRwDuTQT3KwshGucJTQ5hTzhWoF7pvB+0hv
Bjy3dr+S2ZyjelQq9GtoA4lrVb0EmzX5wFx+5vBbGpuj0+UASvb7r76Xa7CPeG3+8yquvUSQDMHn
lqVQXv7O8EbXYgDOcxNM7ZagWXHDImZoTV+w7fjVa+9Vo67EA4BJx5klDJ+P1TLdx4/NNgqmtPWV
A6IsSdsjOYMi6iiqXwcYsYc405LfhQNlYdYUCYqwU4t0FckrxOPWlifp/uPKaBaYStqsRURNhdDz
z0v8/55jYYgcdzyKB3hVkXmPx/qvfv5cukMQVL/RDm9Z+xCx58W/NhkP0rrTI6eYp1HbmiNt3/af
Y7tfJ5n9AW8DMReUNZkCbaIBiApLll7rBpmBciUE/8/lItgVfSRA66GocLz+0fI5YMODt+53ILVU
QGK+ABtElYeALFpg1GW37vTfLebphjKDd7QIJDEZ46nkv41WfBn+9CDb8vWqaqVR1mejHk9adqQT
120YB0ogmOlkY/eyiJdjaf5cBW2WUSs8caolZtMjqtcJnI2yNRgk7hG/BaXArvdJqmKiGW/AX58R
ER1oAYz8Qq2Doc04PpNTsgeKCSigwIh0U9boBSaHAFsO0IWnKsEl7E+J0f3c6EPMoO3S5dkNUOll
bUzj5esYQS5tFVCiBFtq8y7mVqlq9ND9E/qQgRn6E3W7AZYqpq73okvjVOr+2MNQiy+HQGbAHTHc
k6zpwB1kK6Rd5X+OgLt+nbQRe8BkCTU/RKNRz30//TxPX3+DaDtnBD//qE1pdRkzKmtnZv5IefLX
APSyTOz2Nn4FKezo7jhbQE3LxjzV38KSTI78oXpng/N2PwkGgpoUFLTlHXMAkOibYPYj48wV/n2o
aLRglRUpwnjeklKScnp/qPQqt5ypYEhZvK7TmrD+WTF4WYghy8+NF2OsdJMo+pdL3BOF6m2R54c4
A/uaQ4G4zWmC5ArL/SyMDlO4FhmK4RjDWEW/BhcEeeDapSI0kuCocc7ddPneIhBojT36RF1WrvLr
bQGjBBKfiez1wpD7V60swUwY1gdDj1qrNqA0qx8wXJReJ1lkHety8q60KQ+cwFYhCE8JVHXKflEe
wwepHPqjWdVycD3WsbknTjklRd7qtqz43PWaY+1+bO1cJCZIcQpc4TfuOhzmSj0rvUsfGU2RUKID
exOUmmln+IBMUGPvDpRumhNq5/GdV9IVv3RaiBo6kckOccbkPdXoZykFQuU4fv+d3Fg7Ia3WSicq
6nZZHbs1P9cjxTA1b75xSXG8ZIBIAHM73PF37+V3bhgb0y6KOFW4914QUpijbtFTdg/WDDc47ztb
AGTQYCrNsX3cJwqz7KJd3WTmlqXtRFy3i9q7OEjrq1Sq2NRPWuYpYBK3X/1GYrJSZtSS3gdLVI7u
TEDRA8VZQINKtG/MIQfr0vlmL2ErT767p4Nc0Nu4rtF6bdzSBLQKGkpgm12NReNF7JnG0TfBYif9
fOXBsJ50N5Rs2O+tAVMsEDPr3w01dSdY5apMOJf9aIax3NVounFr+ZvQJASuDIWD35nXVCCduDEa
BKrP4+Nq/RxvfuShz1oe+VGPGpl6ICeVihPSXMnX2TzW6t4VQyKXV4YeNzrXMo8DacT1cWqk8FPo
HV8Jfn8j7O+npYr395b+/GPFk2rPuVS4VWQGzetEbapOyvSSMgHZk7fktBOnLidElCB5OtiIfXKX
f8IPNi76NYISuR0h1uS5itxDLepp6JxiW5ZyxHxOKBxaItS9MzPTwJC6zDY4oGGnhXOkJrbPhK8C
oY+FL9uia0cwHL4bG1BXVDFXMOn7HVwP+34GCS/1TLLq1WVyHqcs2RAfOKgedh6sypDjuhe48xV0
WhZnMKblL/sI93sz06geJWglUa/qvsrDSAcjsYCiSoYfNXIe+Yr+2t17c4iIINE0seDNezsWACN8
69blzQI9VJ6UXaom5Tqvx17Hg41quzlMa/VsKDeDfMxjWg9BIrB+uCw74kU7p0jK3I92DEWNYMnx
uj1wd6HdVSmEeY/dGx1587pvZCHwVZ6X1monJYK2UatUSo5ZP+IO8sNE8NrbqEeSNOOelOuKkvIy
wS0mn5OwkWeqz/NfZwpJj1hL24ps++EH4xor/WK6R2vaLrZNGPFQlxiVwT1ohfJs0uukrnsMcORb
mqMRx+hSw37SuxbGhRB6phQiLclTepTS8k0dIyjrkI+N7StMQvxNvVReHxSC2b7eqBiqriIODxDs
8oxPE4MO656S5QHbCddQzDWzM9fqpa3wWE3oGaWX6qV7D/kikSM5/X/VgK064xC+M6pTMl30unWG
Aj/LZqO710fLu7Cj549KfhgWeRiqf2zk7KjQih4Q1HxeKcv6TkQ/sXjre+ekXqd19u9dDMILMQ3C
LGYzusgpUGvAAlpAdAWSEsNjgcP22lbKs9n+czK0Je4j/V9KuGpcPAgVLFnzF0kmSWIHEB9FHZ/y
TawQ2e4uRPgcrifQgrzYf8mqa01KTYkgzS5L539kiSpwATRIWwUok6jAYIgyc9zRyVHSjPzcUrfy
oBeYYh5loVK2wqWV9Eh+QzcTp3nnDb//J/uj9Rb5x/wxWG1W0FT7uxvPoY5iUfnRbTzHPn/N4pdO
yqa9aZ3pGmquqk50K/94FVggnpJ9WhWToKi9tjUJteZBOKl9pW3EYIcALRyhhOxoSsKxyw5HHlKT
UM2ShSbBPNNmx+b8LgfVVty7Oa+bpl9CAQUbxO/b3sfJtmBVA15C7VQGczgZCCJl9pziqjp+wOrb
jMabbAdHmR21K17Xm2gC89LUrE3pn6K17u4qynely2Cv3uar3pZ8oAJD7dy/NXX+2DCEhbVTRY1I
brqzkSrzXWF7daDSbQhf9G18PH+8CXR431r66IhGUaai2/6btMAH80FaR8GebAfXwofTftu71rYe
g3KoZOouG5dPeSoPS5q4ut69a/kmV3ZPXCzYq+t0t9+QIFb322OQjG6openzliCZETyLz6TlU14P
qDlMczDBJq27BDEw/NfYUa90aiVlWnihr4c0Ps+0TkoP4UXeDPdMSNcYTlbYJRlehdjlFWInj08s
z//C8WIHEXkPMQp3o4ucZMbEXTZpi8PKEeq0+p07ZIRKQBfwsJwxXWV1R4WCF44DrHUbDnqTK624
ubStrHvJ1FUAplXdJt44T4yM/02uEo3L0Xuw9mhSdYNACpwur+Sz23jv1luCXvwpBdMlQ6h+L3F5
CLx//WvaaNpk9rUWFGJR8FaQIv5nhdT/bS9cEClFEi0FUg7luwPlpChDGp7Xu0/x5XRV1IyA/Z0F
vDbavkwd/Y/BIWgu2Xi+KSu6QswMTG7lc7znGmZ+l4O6IHfK3His4Pq1BVMJT77A9apDNUcXWjPD
4KwQFjwSm/aQHPreW/VRPGCE5n7PsoYYlq4lHVQrmEMIgATzlkF6OZhL/A0T1EbXEecgvogugOfW
ue3LqTIN+4fmVmig5X73Jr9cRncq3J9e+USDRaiJxGp49Y8j8q5XY4ovRgi4raeyoKjzaGRFnd02
pX20NyKGZZbrvdYWnY+YQ+hcmoEqSA4tFYI5Ogzw+VTjKsjyTo3GdAFK/7vgUU0In9eJJl9FXGhK
QfMBcC666LsGMUJmn3qrObunqQY2EVcQUJBsdcce8JLUuU6Y7Tvb+nuubv5Z79kwaC3JXtyqkWvD
B1VDG0HU+l4mMFrbB8mrR/XNkwQW0iHYxceGaSZbZOFqt84tqBSBe2udhg2PZGfwduvfoY17mZ8Q
Y45410S3ZBtvmcrc4/7E8zQ7qUwixHms9G/vo3BG97KjoDnHwo04Y19qp+1eCCuspAp0AlTL5GdB
KbfKGudoa0lZG0MKGD/aWDLShzu1SHd3wSDNEHh6EpXXzMgdzHaOvBN2MC/Du+Fzo+zYK/u4BI4m
PH62ALxaFlEnFBzuJ/VioQoCYEq6JfOvblPyCMNNCBFqw2L38rH2f0YIKZr5hU4e3sP+F3eANI8R
yO2EANHBAI2j5zMTlEEpfMg+rVGGrQUP/SB2waCHgba0v5+9LhKIMNqwMFVxPkfs23OiV/w66Wv/
W+CcR+jbA/W+0leR3VhwdRFRkYDKxcY0UA5XzDyZpkTQDizVjU1jmd/4ChhmBwRuC9jem769ufJM
R+7k1/QKxU64YPVpg+rDBzShdvzdppxknMGNy7Yr5T93Lw702XHb4W3582I1Q2z9TwUKT/PGskvv
xV5iG92ewl+P+Iuwq17CninDLq2XWhqL+jKub3HuBJzkejhiwXIPCLPIV2H6vcVIt99kmYtUy37f
LIhJkwBz5+JIts+9VIEpx1ejaYddma2/NJBhZrqkUfalTlJ0nQ248WC/USobeko8pxfyNJNICUrf
fXR/fGX+I+lbEagNrcVpGvp0JGdbzt0q0Xr+ozIriDczauHBJVBFY+QlRRd+TmCfLs9Fodmfj6vo
AMo1mYcHLFkO+wpV1t9ub1n/XWQ0GOTKJFrjV17DvseGRhF6PFZnhdM50Z6ztWmgI+CO3DRF8ZPN
Eyq8xI5bax2nn7xMT0y6s5RiG12603uPq4iKujaNaqmv8QkutJKfCd4apmKXfmu141t3KHOc2rw7
jElq0BVKZssFXX8o/Eb7tQgEaVhuO52EIwL8wHaiAyE+UociQSkH71T5sTL+CqHNe8y4K+I0TNvH
wVi2ZZZi8rMJR2ZMemv7dM6OapNjIWWo9yIubnoz68AoMamJn4Y+bQXfhqI2LfXlvhKFt84hWoQ6
6cAsmcc/9Ar2kSyCCNgX6PfXb6Ac6XbzMh5xX2f/DWin7g3zIFdTv0kYz+wl3TiaDkWDnaXRNaUU
PbmqJlPVAICILzptEMw2OA7/xLd3HtEd78hCAWViRRRq+BjGpA5dL3Qal5q+JqRS0MZHgMIY77mG
3sgkGRy6Pnv+ZBzTtghanUzHs8yek7kSFFP1ivULW5fQgt2S5qEiFpB6OKqOGnAADvbjP5HZ2C0G
fpvNPJ4vpOS2pS1oHSCDt5KJq0FMdoI6tQqzZLhD05ke/UawM5czifmsuSsr40PerooY9y7ATR8Y
GxWo5a9y3mc8Qmg0pkAsk7yjYe+Gh4lXLAh/COlyfxJMMoo+jn6NqKUOgyJajBxmuZCvFe2PzoqF
f6oPlTwU9Ws9Di167MkUs3I98I4S1gx+Ge4mSAr5XtR/Qk4g5J5de+1eCH43vUuIu061D+CQeGYw
BNhOfZAusGA/7z6gW6Gje46tEZ4tAq/Y4lzioJCuCsx1eF5BiGMt2wbdborLvwdDgYtZGFOY2er5
v0ullwk7jlw1Uc1lIJajlvWDY6sX9kNDNlONDf0EsHhUE/3FYl2eiW25z+PDo558O7+tzcEmst2Z
mizD7nvOY7QhVEVxBVIU6fopjf88hkH3ae0Vz8CucdU7kYmimaioHo1/mXk8SjcDXVpMFW3vrXQs
YjgKY30RXbuJumHmeQEAlrTYLaBJmyda7hoVsPwSAO/R0F3sJx917FUqNZy39TETd5/qqprauLIC
fg+517gPlXzM6Y6gDUhPERXKAHCZMVMSgmAfIc9iJBkk05TnGwxhWV6xZILR8GLM67QN5BGXd6Qr
Et3yivn84u8gslNFUnp0ahlFA2h7Hg/g8droQWJlc7FZZU3Erj6hj82ngiv3H4b9snvBa48zSKf/
jxfvukAqBUmtJpVMQtXXn/VZofpPhfH3VYGmTZWcAvf/4WGxU9fF2MFghyeDeWKyFzW5Nyv2vxs6
RQ3Se3Q6KSd3tUMVYS3tMBWzmx4e9Wt/HTrIKIjq82GyrfNnuNACXltz2cW/rAYBbVM3fojqY+UK
VZMjMtBNyGwUfQqw7WcZ3+gsrS+SxG2+NJXzalI0S6fUQmXihgcwKNo1XfRzm39zjXrj69w8gusd
svrVNHEIbhslpl30wLrckQ10TR9KPWO1F3f/oay9sAxLU5Mn9LIYG2z2GSCHKcTelIgMV6QGFmMR
r1ZdUfeLSPDAjZf/dhPm8U/gKNjMXJSyIjOzU0JtrtkrQESQnwiy08Tpy5fpe/bmDey4XI83Xr9t
HtX6QIlon21JTsW7vKcfWZMYJJcuamXCFbSaDr/w+b69l2tsmQUZXWlSsr9VZIci+8MjrPsvm6uo
n13suXmoofRR+IDjjo/roWeN3wtnl8h4iIfYr5SAbVN3bJMmddjO7AeGjmJAY5xCoQHSMwAfq1n0
FXoaiWgcVvJCoXSSmnX6gdXu5enKj56mPjTeQKVFbi8urriEtN2aKsN88y+iK19pl3bAFeDoCKgE
5ng22fsZ0nrEm2/8/FCIqOthH3q+4a8Qon04T9Mbvfv7FG32D/axpBwoUZntRRjNx4QvyLihApBX
fEPoHU+KXu6lct7YPf/TS4TJlaQW3WcluceZm47bF3m75Pb93d5gtrgfcIHsb5ltr+oGRNzr9jlT
R3po069XzXlvIdUQG8Ef2lU9pRGhzx1q1PKFpR1ytsug4tD5sbw3JJ62ohMPSH5+6Lkma7sAxtSd
/vgLj/8ymt1WjOc8ZFIwBOIbk23XE+IH3cfnAlwpFyiDl64eUlX7Y7h5NiY48y4wWOda0Q18YW8r
NFfba3XaEca7nbtcjQA7EAS+YA/628zmOp60MCjDWa1IsNOwhB+/igVQkK8cZlRkbopAed65LCd+
IfYlHMwBIXCbILDTabgodCu7/WANGLfb9PDYXh/bXms37jgzL8Szgl7CUcYGKay/PY7XQKc6oJJa
2CCXzVI4o92R8BGyMf128uRI0vUJRnxz+WicYYUBcu+0mdfo83LFanlAhMxk5o6hi18I88EDvRcC
mdFvdMYLOqk3XwAu+scyydBv7u9pqr98Lk+rxCOV6ab1iP0MQ8j8zOgZ3Ov7xfXoeT6XZla3F96D
HfC6fmdKS/eWD1xMDwIXvJyf0gZwMn6cjtNk5+4GSyylR8179Dj24HhGa+wSUZNK5ZCT4H/OMWjS
XAlGqKn53shSl0IfEa/wpb78I70tK0RQWoqpBvXGzR2Mf5nThhs3MIycUKDbYTfFdmA5G5J+El2K
fqlIk8X4gXEkmHhIrlsn/McQZOycAzunc0uKRw+go4IEugC8Hif6oPDfz5kFXAdwrDcFTWi/iEwn
WUkdP9Q/gvd25CLzuL2sxPYboF5Pcr7bNO+B642iHTBaod2WC5gcHcEOYt3/UA44VY0yWWwGoeO1
x9Vz5R7fQyGYmP0jvapzyjcb/IOfN2jwaR38zRNPoQ63+SYrfnoTGBf1zQUDLRvwWW/7GwsaEF6D
Gv5rpnYMdyvdUoMjlx/TYfuFAmp5r9d4WTc3a+pJXDcJVl69X4oJj9sbUXVhkIQZRoEZiHh3l5S+
IQfKf7zIenf3sI3XVDlE7WKbiznYeZo02xwLsDVDFpMRz3efexEmKiiVVJcylEvEnakoGYcMPkBp
89GS0xHg75c5wAQgdJ1wXTGMAOj9RIjlfbuZP6jE/+bsKusVbW02GpEAgrTncxQ2p4L6LH6T61Y1
oDJHLoX8wiOChGnaTYJc42JtBjCjmBhE2NpcbL4O31uaiD+KmUQn7xI/nPhGi+goaLdG5lvG9C6r
teSkfq2o2uQnHzZDaTnj0+sMuAiXIzutnN+qZjJdRbRm/1bPCHxo559d1DYmjhyQmx5vf4f1a1xd
BtHKH78/jvwzVh8bJ5A4u8O/RsDPAaNqkC1ZjkG3dLIbaVcz6weqRctBQI0qq2NKRGlZK+c9LHq9
WGfy0WVv2KOOp7F61UfSnfDIK4VUCdk6QITRIfnEZy/OM5sFLcJWIltB1PAtUunKUW7Z7eyUbRqU
Y5BJIaMob+RxksvfQjbUvUoe4nBqFCUly39fJLWQr5pt1V8TZsbYAkOzFdsgpi+C409F9Z7+lk3y
tGE95+JyzJCZgIodF1Vm3MG2GiaZ6nfcagVcn+pyCgYXjU1b1iwIuwMxoR/LlYH9RQeaTUT8YG+k
2mI5PCj7BPIoAlMsj067KGmzRq9kxwVf0FjG2Yy1s8oarDbRAdO7r/oTpNSD6e/q73XiX3nRnIS0
mvl+jwvf2vhMf8Ak007lQNZhIO1FptTjRA0keECPdoF53tIimlOMlN0EaldrNXf5vSYii5suUEXr
CuWzfYkddJkBHOzq/lLjmGiiTmtnwL+4v91bR+PbP0choTWZ4qFln+OYrc0h26vpxUi2HvUS2M8m
IFUkwnrkyAxCdQVkL33lI3g4QnAhfbg8QVvjsl6aieXBktL6qhbF6TppSHdWI9gJjViELa206qFD
FCyiVDo7E07gQtCiHchuocyGa7y5bSVRw3zXhLX1EvfigFtX8D4893kUzulXvMwsQz0BzOV7vLZ3
Go+fQwLJXpobNfxtJTuk8WWMQWZewOJhtSIFZFlo6qTt3pd9rDWbDLXw7gw7ZEQSnKSwzewsW1x0
aAcmJ5wH5IceIikVPk5jMfZ+ZLAPEzUtSHaHHQXR7lwGq80r0hvacI/VKljmgFIaI/S5kRz1qrgk
b6mBlhay8jcY3jdTngtBfmThom3QQo0HXbO+Gy4kwvEDO4ZAsL37mmEaEa4gbqpr/VxLzDFMI5yI
RgwxRX57ucwA7bDq6IPeOw5c1zsZJABUS/g7Qdh2K6/57QTNMBM5gX24pIIcakXn54E9MaLp6/tq
FhLeFgeyjWQJpgU0Roe6hSQw2Fn1wT6bWkxHpjcBzS/CpLi62UO3i8OB2hogMC1z/XRMSeDp1AS9
TqmpxIFBo4+pWfEQWsZLhJOBdelGCjeKBK63pd6BgUR4deaRAURtOd7bwUJtRpBq0zOgxFpJu/qj
L9pWtp2CyokZD1mrmkDF/pVP5yx3/VLNNegB3ekVWvhF2Z+0EmNy+zGvkclMykXE1DHV+Tf6F8pb
zotLbesrDYPQc9eYvRg5nBk18bJ9891KQ1vkRt5h2NsgeMtkza2qK2hDR+pHxVCWHYrLLEjZ90AR
LiaN0aDbUKfrRq7JC09VifyAPyTbAOgkPFBj6D7SK+Dd10axLpebe5JphufSDrrb165uVXrem9nT
sgRIXiCFGoXWEuTj+KOSTckJzbvvAgNULmsV2P0ToQfX8G72rCQvUdHi+PKmqDhC0cNo+GO15aOe
bP12zdUFmjPTE/CRDIuByvg5aSa2rj2pWfSdfgLpnQT8qKRVUSM50fuo468B8DIGhYwiQl9Mhrpd
3bAX/mseNuqqYsUXAabcAwTdmrLT7uoJwdTmXcKxGGjWk+xKzGQThUDP2Qy+slgC+ht02BMekbnb
GjkW2qMcGEc/7K+FSgaqFK1Kzo4HEBvoizmW1d933cpqonTwqAuUBOQ1mEMsBsIE9s5VArt3yONm
Ic5OshkX89wvntM3dcD7nyHWVF4ygOxcNP+7AVpBVZ51rLImziHJJRbsc0IkbGzAEs6Sl5jqjtGT
takim/ocj8Wkx6YRwxFdWqgHKTioH7ec/1moJcQ/tU6y96S9K4kuzWn7hRXKzHsEeypNhnwf1Pqo
fR3Zfol5d3J49hxOJb5e2Dwm2Qy/mPhvLNoJQ1Pv9j4M6wV6vPAx6IyxsuftY8BhhGYBdqUoWuDc
PDwF9CTBqm60quz94d5r679pjlKvKayaisfRc9S+zmn4kx3xfi8RODrgTJu2sNhphF9lWWMhSzrc
T0SfUXcoF7ky8QZghOF/sSWRpLhCfXYPisbkL80yGi48YlMbYU2VxABLoahOD9Lc6m3nn5ETuc0B
yCIHNxphD0+2hs0UvCGoLNul+QIcnB3nOBoYEDio7Vu7EhIDD8H4v7SghPWQFk40Fe86GHltLx1t
/ByXpQz6rxqZJ4sM74Dp1XzQW55WYeGC9yLWA0sA2YjBLH3RB8W0Jo/GjVRaN0nx8upQQ0e193a7
3X+a9+XR+pBZpBBXDPaYzlsuRkW2SYucHSEUSW9tUln4xPQtOc2FouroGpbDiHa1ybWSiPcOMsGF
4wEMlwrZtMPHHt5zNKOUsorg0818WmF6X0WFTrAjyLDwXe/muX+4WPUrG42yEV0u/kxlLmUfGbHK
4CVgQhml7GjxKaSYIePkEdEyDKbOI0Bq0wJoI2Sg4yDsS/OUH/Rs5qwYZ1/MHnHS7/rpyQBw7KIY
i2fueQqWvP3jUHuSlGtNgUlGuKa38qHee4Pk0e6ZxDadpLoUoDmJklWvXdUVlCPpBGHC28BjIRBr
qKwfmScwv5wEDJMK1dxyET5q1ya6SjNNz8pzEWd/lZ4idXuNF5eUCrxLr/At1YUeSpM0Jy0QOJ+D
IIGip7+L2CDzMXMCyrkw0N4Ym+cFPikkkkZcQT6cbNho2V8iufkT+qhPssvw3jrIdJwvcv19PAJr
CYZvG0hmI/WvMcebJ2AuSe0P+KbfoBgXS5onepzsFP3PnAzA4FEYmZIpBFiadSNnCsFC/aIU6eke
2sHJuVosX630Q2gl39gs5CuhHtU/GsRZ1Yq6ZRgrNWm89/aWuR+u59lV6+OR1yyRw1RKt0XGLWuA
kj+Ja057CO3zH0X01KHp93TMmi1Ws91Ebn9/71YQgYt4XMEXwHmBtbrffqcrRjuHpey2KYYktJcn
N34l/fDSCQraPZHvba+2feBfouN9YA9RSSWvOnIRN1EqsnFidm44c6lpwzZWfHKJ6c5u/4a7eOnT
5/yY+rO9c+TbMB+CcldUuVNDzObSU8ml++pM+NozKWkhllD+MkUJPL+2QKLf0bt8sRi8S0VGtb71
rUJqlmNMgwshO5YXE0SpvXr5WMPQr6lfJqX/fgzo8Wwqnbpe8s9d7Xc9rs4LkQ/IgNbjfeFo87pI
3e+uebY8XY6ZBU9Ye9Q8BQjaHa4dzNsK0f/ZYjrJLepCv2K4U+XDrFuWnSumD1fcfo9VWqDtrKhJ
trhldEfvsDuenm2FlwOiCKARGU0p41jQTxq1elQDdJf1oxlQqJlhy0cwJ7RNZmPFxfa+DIbnojqv
18mZOvE+J4LzcZgKRpX1g9erIMkQ6KZYGrwbWzf/AeDyW3zt/iC0Fi7edoZ54TnbplSsOP8dkQGr
EUr7AsF6aLM2qSMjt5N5LinAgqucU9sfdZiOSjv9UkL0cc9bOwwsuwr6s3WEzWpA9U39DJq5iHzl
CPK7rXaFvwGX0brU/pgqYlA1sqoYQu6dpcYAvW70bJfTyNT3e5LlzayoF7hLGvIva23/EoRPTGGC
M3+gJjwzGTmfr3hkI/PgAodokP6/fxS96Y5pzNxBeu7w1k19qTgwSsy6y5qbeBy5ovAg0hPa+IFA
32RbMxL8APrhxqfnvWb3fMukGWOH8XWDLokYicP66LtlElttQ1+M3pH23SySltwnjChJcisBGsxi
ugTThCGmmyahLWCit1e89FH+wq64zyx2ZrSALAbd8dr6gc1uOy87/uWnqLq7FpZt0F3/UMzjR5Dw
/MBTaAw8OiKPEd5HNPhLf1QvYJ6guq0WivvD1ilJSSNBxIhz2cmzlqxTx0EO8C4+9dJaIKf5n6FU
E/r5CbDqQZUx1EtBLQDYpICppAQU+XtyNpt86/bYeJDpB9Dq+1YULiQEOkHK//orSDn3qOmxnfYa
pFEOBXpHFtB9Yga+ktDcbNqJjORlH3s+rXRkPl0Awzy3IZW1grSwYK3YTkGIpPLnXPj/hopQ/ut/
9qFMx6c1O19gREcnsz1440mx0ZyA32Q3E6YYstCoFjqikkgTSnV0Ba0zGDN7NHzDVp99I/EPTh+B
qrKw0sMvQkPJfoOt7L+A2wKknH7KXrYBDS73GbLo4h3SkRGWxYkcwAETA/o68QpHBSs1PWaafaUx
Q+BMYCo8HASJW4Q5x2vt8OlhRoSjM9BZ0qP1rwu6X55zQpQHBTmHfx1r/136BKaJbKJmC0ulUQNx
TlHpL7d0IZ3b4vE+N3BBb2vQZto3fORAOeQIFPEwoZzY9yuOFKKoGUHHSDDmwpmSensb8p+V+uEn
cc/FX2PCk8jwRUGwmi6r2AgK0Jma+oLmf2ZXlSyGSsgBeU/dy5CjgWnPA8/XBE5Qe0y0Q+tzbJ84
SbkPAgyuNeY4Y4dYCu67BuXryf45+TAVifwnsdrX9Wnz7y+RnhLQo8EZqByeWVf7Q4iAi7WxxXDe
MFtduqRUpyStQ3OggxsHohCdvCEQ9ZN0GiISyrzkW/KWCuGrJ3vCxh0TxlWUO1ugymqSkszzg8rg
1XKd2RG262cE3VD4D1/uP2zmN/XsYhwi8rNY3URkSyeqNeBse9NU477laEFqHHNkSo3PPy+hW+xL
fT8c3eF7AtvzWOOSXIDqKf0TBxguQ0i7n9WSmV1brVNuKyHCcDr3NLerfA4xepWPXCBs1TwfYjfN
UjRQ8nuLootZ9BWk/u3pT1he/sXM1YWjmC23kPHw3r9yS1nwQqu03Gk4B/vSnSRRlx+wPpVrdRU+
RGpxJ2XP5auORG+rhjazFdkTSR1IbqZ6dpyJ+578kzxUWHAC3qKPuKS0/COBBVeiVChO8HsqT6b6
pEpbDeS4lousFsPg3lf+ww7iq1qvLqm7k0CcVYMfV5x2WRoFBVwE36A1FSs+MP/4CHoPiOUN/X3V
/M99a+1vlttx4JTvjmwmoiQL2GmwXZgW95jGkT19f5mecl20uYl2PJmM1B1l8dAVFls/fK7yVdKK
SqDnxI1uDhALeEVnquL58Or7TqIlzgr+qlzuCNeIZIJs+xDMCKTiJkACFBGwHoSB8PQ/wMR9erqK
u44cN6Y/Yq1CYIz9htEWKl4Yg/3488zeRFzWcuda1I04xp70Ozeo01wwZUfQyofdS4JpnAY59e7L
4WG2NleSjwMvx7CjhIzWrhUsVrCJy7VXxWhaSYFQ/r5Vb/J+yRg9WEkkerQXOdyr+9bU4RjcRd04
G2UyVaBs+UZbOSWa+6ub+C8HRTnHznyOow+1G5jajvWA2nNvFTbxehbNlab5BHA0f7u7WYZlPt+A
l1E7oGuW8OTk7EdnNfGbV+mjTYPsk3p9x1eqLtTQYXKukzQ4EhgThUhFIHY8ZBb1iA4Q+vIyx50m
/atjqa7gKqEV482jrqbiuDc7IZRm9vjHxW+MPbnWI1X1SbgJw9ajDe7Uk2cAZIHcWIupK4QAFWdK
ssQW2UXcUqimSb6TU3O72e4EeyP8YuxMYIYCf/sl7/TZ59uW5/k0/41boUj/AW/VR4UNwdtm353X
/P8t0dfLyiaQTcnb8wh4n0bjOUPGqipzppO99Wiz7JOJx+gL6czdzaL8aQWZsXt6lX8DzP9aXSKr
1TMdRjgX9YNhleNwifRWnZUv2s4nfhfbv1HeAiX6Oh2urbZ1MNQw9C4vfm1JgB8yRboquao1c8Cd
9Mo5IrrcmtK/KZl1MDirPhlv0lymoR4Inth1+Ykt0mbi+gc1LfiUdxxxeF/cMjE0u4Yck7K8zAOL
wxHXPLiSNO1kw/kBqiw91+0L0HYpOgkvvGGddZqYP7fS1qJoFQc5mvxAPlU5EYu8GqTkv7CSAZns
F5bzwd2rNOVE2nGQ+rN2g6TCDSHsacafVKUEQPBpP654ZR7C4rDeXYif64DRUWVUguh10OlQr7wQ
S4aIvxrFZmBc6NWqMa8qXpYXUx80F3f25pWT7sg2+YN46VX+/8AVHKiCx8y3wdmsDFcm/LZKQgls
/624YSebhsVdG7/WVu7GIvnZiSgzr+Prj12q1vbn5GaSgs2V/UjDtFMOkFkTkpBbS6v5+mEAkF14
EXDvkL8J5uh6IcdsoVAjHrwcdXZLNENxzVM+vT3mSNL2NzIcK4QRrvtFTCvFKYMH93br2oEx2ayd
1ZPXwqyC/B9JVJwChS6CZAUcrEcTlmY6rDIfFegBXDomahG0WI2Ma4uR/7YE2AN+wE+YVSenDQIM
MYk5vIq90rJze8smKsssOSfrlr4O+4qUAIljRa6LDgj4y1u52xT6vvmn+4hIgQ4F0WuZyBeq3iC5
dKq74/d0rjxmVTY/Je1eaMBXH0n2VKYIuOZVsNUZuET16Dk4lOHN++c5MFst7h4XFpltp9IvtteI
03HSqzmcpuJUWiwMtWFV1tkAdVETmhYIjx6yFCfW488EGDwrhJi+5ppxw4FUKCZ4b7tIiJyBq3Y5
LmfByCOZcD8kmWTD1Y2xKICYJEY4zvU3O936vDsNoeugqfiyKiBuxhu2uyurgQQ/ry3Noc/gS6JM
pseVDuTp29WGarBexW2b6umFSRqdiq1FZJo3s7rSRmbaq+knDO/y75YRueHUU8h8dnFRsEV+MkWE
N4NSELSC9SPInzHyCyMh+4gdCH1onR5rVP7H90mujvbqU4aTILAxPMnlxhnx5bUuJrLTThD87QRg
LZX7kdc39IdWihfL2+CV2liw+IAisRZ2PFp0baMyLHC+tNYYHLlSiBCl7qqQaTkDVdrKLHh1F8tq
985AUeVvAIoCt20KWKF+EpKIcAuSNfyY5nnAG4/fXuyHAErsLnO9vdVEpNglNm8XENWVavtTrvn6
vvyFODuaWD1kcSDdsnq4oxigMrKXLpa5atMy88ZGwrYcgUdc537GXoL7VsvdA9lR/tRYh1hTHgeS
U3zGzceeVB2eZP49STfel6EbHWU6tZLqq1G1RFIsvA2xb1r3YDrxPkTDFAIbSnk4uO9gv4ryt6Dy
IL727xM0Xt322LDgq5C3lZP3jQC2RRnRKl3soya5gQLdcQQEK/4Ai5vFTu5iqxsML/hApDhajlTq
TWy7w5juG1dGG1hFAj7x6YBgX9a70odfB4fgeJNHuMc/466gSKFqEZ39eHJXkcf70gD4BjiwiumB
IH41QmgrmiHOmNqFrO7eG5aYptMDzaYv+1hpjTYnyMbylKc4RVUkacP96bfCxDnHVJNrFjGrXh3c
bWba1c+54F3k6CTwEa1Gc3mwWagNaXg6/w3z5KCRh6dEzqDsAoK+iKEEZOeDs3O3kUAHW4jZxmy8
GPAMVUEWI1JRSkfC3s+7FBzi2CGMGKBVuIa7lIcGc2jjsjJ2anTPbpWYGXvkEMZG2EOwd8NvHXQc
wya57Oxte7bAaX7x4+Hguw9fc3KVSvzXK0kJNWqholqFfyeRllQh/QH+rIeedsMOZtDHl0QRvXpR
2OGpS9+AKCNHGgYJ2qXkXV9ED0ZRHST3/3wxkL1uEzysdM+rOtwa4MFyMs5fVoc83NlsiPpKNYPO
yEFsBUtmVvTK3zo5zQWrbeUAUy7gc7BqQNAEGBYavDva61FP/usPFO5FRXxNc1xptjjAqHJmsHoH
jfrErq3NI0Hv1Pblnu/Jgm/gDImfZLvYpggLdK4CYeIYg35sKs+PNkcUYcsjQBddwladiGZD+KX6
TFjbb7cl5zy/TcY34e7AD4k79kY90A6A+z4r7YyBSzr029Oeet9FWRSrjZojHVGxX7oPG401jUNj
c+PA14jpeNUNh+PPH9/81flrxWKltJLww9p7KbJbjZFMn8NVskkUlIj1oAIRTk7VO8agaqAJFutE
0vbVvFLvzjDRJ5xG4NTOBXu+t8bA3voYAgdrSGeAmQ3s4s3JBHMwQlNag1KzMhMTpyrniB13Pmvb
kgQFkE9NjkFgEVTarpH75kbul/WqmZrvGwem5SZj583XWomfmNZ7PcHahx83YGBSSX5TJEqpM46z
uqNup1medWD8i+WqPq9r00fKSn74hoP6ncQBG49npxhFkmn3N9Vylr/Alr82H9eQcJWH7EuRoGHF
ybM03ghqcGJKi96DLzKX2wFKBgSfoG1o7vCN0tHrfM5uuWqF3GnstxITwpTqThr7UgWwMY4jDoSB
83f7NtZq60Du88EplKOQaklNG3BCi4BneOkJF4hY50xHzPajOyLQ2OceBHWFiCQCxs6xvrWubMvQ
YtykQcTtT2h8scfsfILiJ5QGmaZFPrZLdIajQZibWXbRAxhVVtiFTxACfH4g9HAOq5rlTofUCk3e
rEQaNGwuuk6PQnd3c5Z7WbxD/gPeszdrKVWYM328TADFPYhg78h9ZKPZQhKmHof5Y6keaI/ZZ9W5
zo2DTSAh344KAHaUdVb47nbNciH4jgPZjr/A6ILRp8n3/4ACZLhhnK6fqao59QYf1Jnxr2Dh3CNE
MYdlKYNXL4m67sV6Q8mizU9P+RIYEN8sVadUTYMmgilJ8J1KiAzaSLeLBccAp+Ch9SA3WuM2nnRG
ehw+C/73qnQC4Fky9OPDvF4Ym6Rf93kzREFkMtSdhTMCwUSeHmOx7gzZpop3+Ap+ASjumhynplFl
dL87a9IVpd9fyNFTxZAosfE4e36nNankdhlohBskMtSe/R8c0oKtUF0BmRXonPBU4LXzQLYuPsgk
8KfHtuz3aGchN/e4+HosJe01wtcAqsxOycjetgOFo68lsfaC2ox6RlpDXpfyu20kZeLulsYeI0Ai
29LLIcDDusWgeg75W1yLdmrf/Aqh5aYnzZdmiYVB0680LMkWUgLtKaqS8G++uRZZGEif/vlrxrLK
f3V2vlmZMpMcPSiD3Ma2UcCWbYCv78p6r1ylweRaSzodd7lQJMd+BEQPgdGqfuTy5Rh3aL9VSk7E
6lnrEkoWu4HPpNSg4sw4HfRigooc+5pGLq/0TgH3YB6XYbxUynza86eTU+y98s3t0LPbShNih328
OUWeBNgdYLQCs+tg/+djnJmpWp2sv0tCVzKUoX6cFdSGbnWas53e8ZlCNOxM2EPRKs5xiv3PotkP
nZz2yjUv90u3mfWGMUppRdOwH+udXA9aqItDnEmUl8CIBOnmZ9p2/Pj+6UtN/mugBpe86GvbyHwQ
aV8qioSjg10sx+VXrKyXm9xIbv7CqJ0d4JSO0YUq525F7iKUtZOKbwy4JEOiRDJIKpOohEd4ZMQk
cHeOmPTxzeElBV0FMUV1l/iTX+W97MupxBR5KQ8atYZ37+kPmzxFQDBxvlKiXSqTrjuSpjfTaxG8
nk1GThh8L577X0QoanUqoMnn4yEx7qhxMM9qlFHXV4y5aJqQZdKjx4fc0s7xsOcqRoD1RVSlwZZ4
CrMSbVS1UKr5wXe9TvKfXX8mcV0I9wp+kMr/Su/OLpxLGLRt4exQZ/BJkVfw7vinhNFud7isu3ai
4LoHuzcj0CO5FnqF6zEERWWL1i7+sGrDroTudgxq5qfH+z7SIACzgDuHKl2o+OYRrmCnzYAU4HwA
bMlHgSF/QRwZBcnmuCmZutkDFi9y/b19TTtEXuP3QK1HIMNnz62GCJKpNh4Ioa0tnH0PyGqm5obd
i0hbGTYktKUflP9WjyfNx30dZZJ9uzlYXMytFwiivzDNMHh8Agdvnj6jNLtKcUX8fwbMxEXbBFOX
5S+/uhNIlp1PaflNFKRqg230gCaiCx99vTSNpgBogibycSZUKefwDZSfNurA45NQQQa8a/tbaUfe
EhEIH2tSeqbpQoyCBfQn3u/PTMroyv0xEnePZ6mXUAwabY2zBohJ4Zy04CfBSVAIV27pzSorbcU8
vw+qsxM3shsUjZBaZINrHS4fbaXZ2MlLJMjo77kVqnL/h3RL4ROuQ5ruvMs6r1q9imTsN/s2t6sd
p90u3SBgsqk82LMXMRlmE4/U8vA859Zzxelk9X1N8Cwwi6BvOVv3u3MYJqaTmozOY6sin/KNkItE
BJSWoMZjvMjpSp2ghETGo6C+jfHg3Y0p0u/DANF76QtdgVApl2XNTsfPNUrRvn9hiepgR20h/V+0
/MDjbcUd2k87MRPwD9O6ZUJYwjU8vNozIjvEcyKjaRoZUbVsmnMgiJ3MIxxz6DNXQLKZNJ10N2Cv
pGNskXIWtqTMs1usv2ewVf3hs5u9zZLd9BA22UkDShGsgDtml276U/6ha7bKyc2ZgA3xkEh6VO9B
dRxgCFcfk2xRLxHY7sNBwneEL+u6m76Xu9n40kU8PbwH7Htw/aMlgNOyN1hdE1XPtVL3bJMIjukh
US2FUFVural2+TNMVH7QR/8MTG+OiL2s05AiIwlU3G6hOYoK9E6YHFvcqw59zZxJvNRJnXaPW+0x
q0OqTCZJ7PNwBCg6PuAZ7g8uAZA8cBnpZSL3liDcK2SZ18peCXBPzDv0wwFuxkXEwM72O4RwL4h+
pP2uslGODQh8YikSsPAXUP3cqGnnTnoCYTr+zfJLBzSR2rTvEkb+ALqyFnnYyhFmGTWoAuOpixlH
QYsGREylywBU9RUIGAMEyPZYFEjg3tXY9uegjYkC+wSN0Co4YYS6HG5CL837RD8BQ+kCaISGrYKv
GfMoxRyRxSGBvuD2Sx7rKMknveKnFuoHTghmHdGAHt1YX5J9tgCmZNkXMAlhSGsYWJLE+qeJsnRI
Uv5/tSuB0dRuDhuOR+XmluDCJgVETdyoHlR85Mh5Y4+R+8SV8u7EHaqZls3nK9eKIhvZPjRLMkgs
jfQKJyH17ibXc6EPawjKw1sZaWFZSGNCQuQTlYj9Y667lWpBbVurlPtdr29YEUI8wSpF34lvqrVv
IKzM2N3hj1pRTQ5Zk5rzgX4QDkxRYrY7v8YWTrTyXs+gwcEWet2ftkAiC+azgbXr2fJRfCALxy9E
74grS2IOJIbM3QtGBM1rHNv4dT6CYAcyrf2NuFiWoidYfnI1ckrmB8Hoqzg2nxd2ydOPTV7V1lmX
qU9lMHib+Cn8/HYNVAc1wgObtpJc8fqpM5b0txiU+G+05neimbxqnZsnB+Qd+JkJmneB1b98Vdmh
5T9HRgXSKQjiKqVvkxu9hVQWjVxKeQoaD0vboFzjsoR4VM5GplwZ+1qdOwvmG/sMs44jycbR995v
sqozvRkFTASqt5J1y+iWou3E99a8+d28AqxYuo52uwXpvfTQfYu/ekG3B4dDQFUxRG0EtsHoivu+
oh8GCYbZWzKNvp884Uh+NeA3TEWr68JGQ5LRnjGMdvSk1tD/U1oJ+Uxy92uXiZSuTfhFNqC1lIJT
F4JjJeFVo76XTe1J1WERbWccXmuSaN6Nj06Vk+3edsNDZYIZMYADeM8LK+qF84qpfhYz3VJ+vXZB
OA+zoioCenh4DtNshr2COIJaTWyFEbYF5t70RYw7fQDm8UIeCHM4Kah9kny9koLz1iR97XOE4pxp
SmSW8cVXPxfQNnCE8vIhEcM40a2WYwVjEMTdiez93PsI3zZURpNDGGQakUMrX7uNxXUSjg/TmzS9
GNfkJ8xa0vbR8bjvqzIoHFbmA75rZo1Gb/jUzerWumuxVp+QFmOWVWKPsW6sGToMVbXOgpTdwGyP
4ok0sjmfYLBd3ZxkC/5ZkgJwDPb2dV1GkQHwpLfs7YwMZkUC6WCV45BUwxwHJoNO4ay/GFRc05X7
iYnltJVPbXZYJmLzBURf7pJWdFBs2330aoXooKET0CuFMC5eo3dV0DXekweDWlYCqYjTEJeQQohK
5RxHNFxWGZ+JLH98eTKNRgU0ATJZ2ZWwn3dfm8fPuu6tqAQ9C2ynSCy7cSgCBaqzJe0RgafXZHGA
0831GC8Qp3f4ogH2W4K4q8VTKPfHXyAa4nwU8juugiENuKzoWWZkQnV0Lun4MZP8FJvbj0s+OvVk
Boyzc6elveLX8Kv3HfwLqzGZSE9VhMsDHQ9eLPIgC67Mug86E04AlulSg5MD7RPb2h5yMrQzTIr3
BToysoScsEFxr98YWwtSaXAusw6tuhJusRwYok/3tTmlDpxfrWbB09xvv24+xI0/ZK8FwqlbI5KN
8oUN1+oL7QSPnBp2XbfIE1lcsFUuOYtTs5/UjXb+YxkluNf7J/S6U6mwCTrImpV4vk90llVtIzGj
BiFNxEwVLp97yS4Z5MSfbUqVeXKGcInMaTls6kGJ96f//N08mF/Tf23dUjyuS8cmvXLvSqnfgIpp
i9mqq3vZzbb5xwNVUSmznE2xCGjMzQqzTh7z8o8rMX2PRD8koWa/ugKIK4WKurEyKmP7OL+Pb6N5
QZl6QJBiJdBVN+KojowJOSD3NogrI84OvVUr9Qc8+D7GF7JOCQiGN2rdJ2qd4U5/PnoAHwN/qQlJ
vpiNA279D+pc0ZyLWLs2OwxrEw2vAiZ391CAAXFTXR0AQ1aEI8kULtgMghwz7N6wsbo7BsbvTeKU
ZnO3gbYf3ug7O7zlZf+5OHkMWa7R3ib9WnHpvr9BLpnjqYIUeulbagRb6EhRmE+rhYvUllm7fkxm
adKfjMiWwEXKTACYr2ZEUL2js93GnKkkSrIFpi7184h0wr20oBKoXqJRT25zOMOXisFy7UDDibOE
MQio5uMyyKUwwI8Zd2CM3wIzqZrYcEl6L3t0jTuz8NKyd71eZKqTD5vy255o9ygRl1iWl1jxV+LL
gbcFWSKO4KgdOu8dqZjc9j0+yN7jmHRmlfWqTzmk9ENL76269f+Vo8maOxGRFtYujXOGnk32Z9Af
6fzlJGe546iOE9zeopC5taiNSPXUHB+W3kN6/UxCxPVylfWcTFE3Wt6OMHLHqrvKPWb4rCGs1ZvK
mYQHioGyvqIiWPXgBNLpBV0ZaMeLQMkxQgwUS2z9e9w9SFRwNYEEE8eDZn/eUcmv9bH5FLZajt3r
ZI272Q7bRxUpDHWrmm1BNQKU8atZnhr6Gzi4lTCEGsIIxouVp2wu1h0d99Ky0IHl4Hzt2hxIEhAS
wptnspdZEF4Wx5tWDELYfEyTtFUXhAnE+h77m8TbG7oz3bbLEtH168VTAPf2BsOdd4JqlY6VcO/P
M35qeykNcLD9i8E3D9Ag9opkWW6eJYmsH5difhYBPyuZ6kSymvyGTLe8W89dZWzzKnpN9V+6bGV0
GIUxYqIRI1Q5TRNK7hM+KaAtT89goFwtyyDfL5OKURuhzMb8KV8z/yMBcz24qbVNpr/HAe1P4h84
uwjIOZb6/JfP8WJXAUNhr8YMaphlAEbQjjh/4hjGh+Nb1Mj2991hEE6IZBTRfNsgMOBrvO6SoR4U
dxESqZNwnDYJtF5QwYJUKo175Gix2YmWU6RTf4Q4yRbeP3fA6+8oJv75SZO0SqyshnFcZw9HcQKm
Ev8da4cgIlu8ue3vAFQD8qoNk/ltxl0uxXGotCYR6Wdv7TLH5IgXIkrf+VHsRLlQXQaiz/P1Vail
w5m2YMpRhFYv+97Bs7H7lNPh97qG4cYahTCyr7DrDYe7U8D6qWnsJ2OGVq1g6czsPAnTYktrOKnk
vN87eERU4O7E8eH7u7HNsDCj7T7Z91JCS+Ieao6FYu3GENpkS5hWQVKpEZXwhxu7V1a2/FrIa44f
o9KziKCFWwkvDkRa6+64YuiN2XPTxWtX1Qj8Och1HfBcjG1y5soOg7qYoiHOmKcqXl+XfFQLdr2O
YMPXtwbqQrLrHWBJRAZYM0Va2Twf17kK1oh6aHmlEjYpILxsAd20ciezu2Ssx+/hRcfwBqZKluni
Aeg30c83S80NyyBQNPi6A7PUG1RXqK4NmyjULr/qSrirNOs/OPEeww8w6sQN/5EGWAx5re/NQ3Np
w+63SX+xf3MuSxnbmDXY1Azhim2sMfnwpbVUhKTIgkWe2MGCQMOO4tAi7noxp/Yg5NcenuqKPrsu
UqSdy9ihD6u038YErh35nSg/zLEM6NVgvAcwPHS7kHbM0BH3CaZxQ/NJfRT0DujF5siGKoaZJ5zv
puhgsZddL+nXHxL7aUq1onepgBwTd+OJrmcRPrBchr6RCFq46h1GaMTnGHjjkAes3NTlZ0NcssGS
K3qJUu0Fh8To7cCOZUkxNZjZUgJetdA6GplrY070AQr8k7HSC2o4a6pwrr1HMoLuQSGrn21Msq0q
IT/5XPd11riOhUebdKq8ctGGQynLdrPUs+9YhY13J/GCIuJjqbBihXF83OYPXzmgx9Yv5GyxzD/A
3r0etY4rWx4A/YxWzkUNzrFtAvgqkdtYUobmZpg5+ozWGjy/w39RGPTXsNFK5la+YAoBVCJjCnmp
RgPgQumJVq07vCUS/x/51mRaIPsFb8OeYkHFj0DUMzn0beLySaoIvuMsqP/IHe7jeVL6DHWnbKdW
6djo9eUdtontJXUMBRjzRIOSwMAmKnfIR2DLX3T9hAmMAPEGA/7VUMVHUz/dyo8gX7OlXiCxGmcl
8Kz0Qd0Uo3GWe3NYDvEV5hLSTmnUeEIzqspnObK+wZ5SRFsz4gLRt+yAgpPnGXtx8wejtA6h2U8Q
wbr0coLmTspX4ujRshst2C9LwARsrIjSnDV5AjGPVHyYe3QUCEoXhGi/mYwvrS14ACecXWMwSP8x
BIdMNhf/o7PUDUSJO+E5oDA3Kg/XKaup+BQ+eAxNRz6BeWhMb08zkb6uoCmQZ3rJcoZcRaorJ0QN
WUtHowPOjZtUVDzARFIz1mZotJaFSdnfiBZqRG4hkcJEFiwGR/buW7TkOsHnOd92o6LoS9yFw1jH
u/MXiliuCzW1H8LUHML+fvY0Ms9fG0Ng9xFYiqf8zLDPh17n7JmGCmjES8sof7gDygl7QrcIUad1
u7Xa2HOlUQf9ayE7aQ2Hft6nq2cXiTKSpR2UPdBUbkVm5wKtOidpxokFWHS8CounqKbCYgjcb/4d
vrhxgW7AP/0Ul92LWeLtiy/7/GTX/qqNpvJdO6OckgaLMiEg3RcdLnxXn05nBEVY/QqdorN8lCYT
yaVX5OBqBHybOqH2qcRX4llBBgt3lOpVycae6R7H2mgyI4faHRo/Y9IRxa+/b6MR6iAquY0cXq/Q
VvSSWih4tJsEUcrNKBU/ghvmLcxx2CRylaR5Ne9qrXq4152jJJyNXNOv6LuT/+PTwOVdxy2e+yOJ
VuZi3lLNTYrl51EvotFHTpg83RKqo5OGJYN3DgUlYWWHDQy9YGZLfBVIC1M7yjbFrlQz0Ziwnyod
SHO/rNhCIcLAzXVmAUE++YIVnPtq9Y5vB6R4B4++3ejsmqZdJEIx4SNq92rC2I9e2zVO7flhqIDK
BxiHWbebauHsLUhLxqnpBqbvyu1ITF2cMk6w07TubsITiBIh8aXg2dHInT2PPz8CPxQYY/113uxC
SctubF/xnx35TbSrqipHyo5v6/fAxa0aRBBtK2d7URk7fF0ny++bh71L0qBv+R0c4J9S8yrE3NFY
lrxnWuVWJqlsklyFPjDA2CKvXPjEot6z86Yo+Ac/wsvUs8r94+GggXjaqMvxLXD4e9mOFoWJm62T
1bJKZx0O9sbfnWjuSUw6MKs14/49nJA4X5HD4PFtiQ258e3vLAbSv0xoYtfw9/eG9iaEm5N1auWQ
uf9ivEfcXBOaYWaLlf9x9cPDsxaMfr99DZYON71A7GVXT8jCNLFqZp86CpANGUzeNy17U5CNEC/v
CTluio+gyfb7NLBnRfjjZwPwK8yJC/a0BnBEFAiX1CCSavn/0/ErWxRpDOmiFnm6RitjslqcdJs1
TCjCCGi9T74DDUWK81x2gGZoNe7OkYxanqwMK58wgKfqDMzsuCpXxQieoZCwdDWzPe2pzZ7IsFkV
2A3xcYykmngLtjKSV/WNirnpb+r76XIPSAy5zgbaQxd9mMICyuAOl36cHKSctKqnJjzDTlNpymNM
7yJpH1rLzTgNkQOe1cTNNWAA2a/MyuL673kk2Pu/awqnSNesOMJTOWHUtzcH0jwa6xrACMzsrRDU
+IA2GfWhp43gahrp9KmNo4Vd6hDaIOl34lRKxiUlVxWGROivalbLOL+HmN3gwEVVJt1zfeS0t6rU
oZciwT0uUJFZxDGQw58IQFyWP0aXDdiHTEn4/Z8kzMDXVZRRljRyGPmeKyk13D3ZEnbWb9MLSouU
LMkJTwwHd13t0MvCHrNQcwzulMrYROW+2ypiXrRpxmKjGSPH9QpTa3kQXiH5Xn4epBv/IYP1RU22
Se3dI6fAw7Yp/jzb4t7fOCfsSEmTwQCJr1wLLzSx+7h4y1uIN6dUUdeUXkk2hS/2delclwyMCmBH
E/k3aPyI3luduTpMZn4tpRHNEgQOD1nWCqXn0TKfuqbULzEN+o3oD4wd5P9fgkof1CTBKfWblcMR
cYxinGE+mkUrnrXW7VvNwgwL60M62aitsIzKiTXYL59lJNQqm9rUeyPu81sxKompQU3ey8+pnEiV
H/vslrRD2IBeuEkOIQKn9G44E2QER7Vpo2gD8TGWkz7YgB/oyNkTAuqm9lC8tUZfDeo657h6Bltd
clkIAf380eu32G9vq/bz8/dVLL0jtq3R4orwUHxjtnCKqHE3BEn5gVAKRVQZBJkY7aWhxQL52Yja
owfs0YUXS965tjUrDhXrQNQjAN/JcnYmfytSRwfkomTzv1n2DLpbPPGfVhjrAHtZU5i7NccNskGE
j8AN8uv3xkuyo0Y/LMMCmm12EcRgpNtskBX5dIZXi/zCzN5T4W8fWYQfyicJEIqEFXnGfIwWLi9a
i2PVlkim8gXhSWSFgATRQeqTehQW+/aKomSkjAhMn2sjBQmhPfJ8SvdCt060hX8pYSj3IW8dt4Ou
0d/ylor+LinpNsrgTMUOosKqCIHU43/x9BDUFiklUUtmbVB2c8GMshhIUdWtVrhHj8dOj19V4Bl/
kvZJQWnBlx+Nm7e35XTDlk83T3r81wYAOgBkw5ka0PnmijDeRibh4Lnbnr6OSdgF2a0JyM6DHwxu
Vzhwfbfl5umRQmtlqTp528oP5vx3DTlhpobAFVGVyv3GFQ1KxdQN8iJ0kUgOrYehHWfsoC1GWagj
0EEWs538Lj/FMlvA8h6NaeZ+p5m8/VjZGu2vTsBahnPDmun6WoSlUfZNFYDUPptpbqTOqXjdtCBD
GtY+OR1HcBLDNnUiA6FNR41vtA9IDykW6yAUFFx4BevTF1cAOkYTEd0cVJApQXc7Ddyqp3YkWt2h
C2bpsDqh0lSu4nR3Fah0OdyCgm3py81l+h9gvJHvScoWWqub2e1r3FfNmEXAcyDiekFfpNPMPz8n
j5QUma/qt7GLPgDac5nl/UMTY3J8bLkvcTlXfhVbfcdYL4q048kARMSRidBixAOWBvsLgX6gGZcL
WuWp2psedqZ+rC5rAiAru+syUSG30h7EP1IBqWAWQJBw2MvQR1RYhGrx1yX0+EWA7kIqWGtN4NIQ
mycv6uoGG1sMrNvklD9/dKfPaWdqTm9ziHdbQXgjnlk4FlT8yIAZ/JND2c+Pqj+d7XKzCFUT1c95
pixYDpeO2XlhBk1PviqPM9usL8eM8MCP8VGJUqzAG/UTeYp1KpD7x8jINj3h/Cg6wXpBIkEorrVe
KH1IK9K92vfUaxE+RHJinK+LPGZodMbGW9Yx0Ifve6PxLp2Uw4B24Z2BswMzGksbhWI47O/OT2Be
lul9Kq3ZdSQqm8XPi+bASbetwVzzTppQCY3fDrgfLgoZAHYqKSK3G5a8uNirBQSc2woEOlliLpB5
TzxAEoxAdB54lHS0/mPcwpIrJjOyolHK2F1uMYOdNPMfcru0NgnDPKAWfBeRDUEoj9c/UWy1Z3ZU
BcJNjRsns//vpBh21I56OovxyyC+gYBY2m+4sbN7g569ExeKqE+RQtOk9GxuBkOI47WrLCJJhcrI
2VFit2+bK50+GMjn9EaZb6Z0uREg0tpREqefunrLyKI894KWBFW6pCBYPQ6YKI9WIUzINhHdoYQ+
Pe4h22NtyR86tlEwJAzki4X8W9BQ8cnpIlPQi+0JXo+y9aBSOm1/ICCR0wrDBCMG7e3TImdGEg2i
tsx8CRwaWj9Si7/yXPkTlf7nENvNf3GqzIM/2SPmUx/Xsc7nMhWCA2XsvI1A/XA+9YBpZinJSvYF
6IMOCNMXym21pBtDhL/UY348RM48Sfvmr49nP0ugryNaf0b/Roq625KXXz0qW13vo4iG1sQrxpT9
c7cNMgQf/mYINtEUAxKlvFF4jcOlXS/OiQbVTbftdBp2/fNl6eSxZeofySTa5ic/AMlMnzlx73ss
j6ChtllKxUrA//nf8hwfc9QdehuuSGp5bAZ0kAzKPSiRQsqm77P+CKNgpGWxFzMhAI3DPeiSmCN2
hcJCkpAPQNoYlhBRIq82QY77+izE785/Ga+FQud1IHZ/WUoG3qck/17s/iyXXODtIqyswqDPEMSo
hrSzs//yoetFg70tv2f3TF+Ky1i31ByypEHL3CuPSmkOuRv0acEb3cw9mE3zdyiOYpyV2DzmO8nG
4ERtw7t5BRlz9Jg/10K+/DdOzk7KPz0GRaPWHHGpgm8b3QeSG4ySMhHJespDGK4LJZgPLPC2Zmfl
5FDk12OSe+LMw7ABsiou7TgBQ1kcxdd7TIuTz5jFvjhGvWQeVYUbxJTKJszVfjLlrx4DO2sdNc3x
9yM6/DiSB0DxfWGK53Yib7Nt8x9YkEit1vZgI96Uw7p0Mi7eFDcmlMjuHLF/OBDYkHAkGIdl/DrE
YWvgurFi7nuG8lgsK/NpePhNyO2dyngHvhnufCssGx9FQT5p1MetKMitunSo9PGsyGBDA8xgwtvg
XeMLMsnsUgpVc28Fpnmi32yF2h0u6063YOv2xkKYsDWmrya6P95ScH1i3qULZe5Az65jUCcyn7lt
1nJ86YWmiJ7VXQ6B8Gou6/rz6Du1khAbC9Hv36XHdRigQ31cINOcRJH9jyN6LGR9bAQws7qh1Fu1
OOFpdKSOVrMq/iSlKXtb44UF2kEr9nY8Q4NJ+BrTUYIp/pVx2TehSyHvE88oq0k9jq2/y6hIizu/
XTai2YHjMLeTTBRZzFxh/6yiCyqVhoJgqAiUD3xWRZUCef/TNxw8zgcEMc3bWN325P7p3/WJ2wQv
YffO5RlTHNx0YKbPSsqSdm0XExM1TSn+v+O/KfJaAQCl0EWFtBN/p8vWx19jH73VnaMTSwLHVUph
mDEliKjmL6hoYYCIbtjKoLxm+Il5fHaX3uHMgCoRavjEevtFqLJNTXfHdzUkmZNiOanbZfl6y0Wj
KjpC2kjO5uPKPFl6qZeLOBZTwuZt1MeHKftYsHi+zBgfd71GKD7R/6GUFPUAlqCtybPN2BtwmRqG
IqgR2pHZizduK0D8waND7O/MQmt4xmOkieVvYI4G9FnzeAVqM74xtqPxdkbCTEqUgQKw977YsRU4
drunnWIO8r4W3EKspA9FGDf/x89Oc7Uyq0ckNCrUuM3uXY0mnjoXVZUAGGSfI93Oclusrzo373+M
3lTj6ctWcKDmzVlv7iJoOUUHH0pvGtCuIW2sj981pZDGHdNBK6yjVgae1IqKVHnduPZEA202/2Nm
3mA25XxFYd9wWDuToY+hrTOPRBQV8rtSXiugDAGGbsfsT+JvmyYitmNPHSkFFh/Dh7YlCnSD+2W6
E2SEnOt2CaaGtbVD+gwMz6xfXY0zarNaswekKmIANl3sVRywD3FHozIVRLaFXP0LMRXIt2oQ7zAZ
l8hfw9UtWoAsOV9RH9iLyAc64NTEo7C/mnA0yDzawwdAZ9ObRxLx+8vbxsAf+iq1XSQ9zYAGkbTI
WWE29nTpOO26CKs95VMxBTf1prZ/G6p52katuR0ORkkkGopUrowKKuHU1GAjs2/39Pobz3H88Grm
WLowXXYGVyWvCIPxATVg1vRjRGFTw7HecJBFpq1LUuor6zFVg2bBCq/x/uP+gSCOzcbkWMI1TKB5
f0qAje9X/qTQv0LURNHfQyid0C4/ksnyqKQAQyRUKB4yHNeKSm00wBZInV05cqss2YcNpF9zgj8J
Mlea3hVK2Y6UtQ9Eqmczxbo/0HnMnlcAO3pN/L/Y9fhacmC3qKguPl67yDPqRxR5st3690fIMlKI
wgz43YpVeO1UYYViy8vOAEsWhgUfNgkk60wbUEX1EyKGJ62nMxAMltAe8kD+yg/ZuTbq2UEZnJTx
kEKCAvY2Yw1CXvnVzq0cjHZjczWzY0PnlY908WBcKoRbIDBH69stEmJ9TDyxkHaRFn0QsZJJrHYx
t9QDCzwuNDI4g3iOl+ZaxpJTNe20lJFx/ETg2yQezabcn61ehhk8BoX6XNqCZsPFSmdyXUuVxPEr
6ziSnUizeXdWX1+jN6F1pAzWyNKkOQrtCvEhs5aW/eC3VDLuiRuoKflJCKQy2Lf9KvtV3d+p4gQM
oNaR7FihKcUHsiHWdvphBpcqvIu/QytOjK4rU2WwwhXZ+mtqRGNvN08qCwOedmMLk7+9NqHKbzqa
PpdO7liqcDhcd8+YRDpWFlNe7aauhYqddDaUjCF9fQc0ZcFxs1snm05XVb/HK3WdVX+rPRl2iYv6
CSM49jma0buKBOqZBF+x6owjUDYzoqtgf2ee15aHOu10zVJkqYQVeEiQwrwsGxQiAI6d+9XNrSyH
MgkBdEA62RADvDbafsdLUda5q6JdCyj8MGgdyGSlxURDpyKH1yila4aJSd3FSbhbVlXRCh8d/HZe
ZUGFLEe4XpTIaIuklhiCi90wyMttCovtQx6JzrY0nKX6uPKI5Sf14DcGhXtYKJzjAc1QSXGrsxX7
3PVIp0DxG1Nz9w4GQdTca9WT4GbcnU01UWhghKnTwNLB5y4AQv4CVOD5KX7Anxcr8trhHwzrUa6y
8eO/6xPeG1n9/FhYCO9EUI8KRUh97wDS2pP+Vu+FhDQJDPMPfoJR/pvh/iOklezB5OR5u9/ri+1G
4/fpPdDN4mYqGxHJ9gBjJ8lSwtRe7yOy3DbJJfQSZKlbnBSvpHh/eNifzPFTRQw8sZ05QDNEbdrX
qyfrxLCo7Fkx5GC2S9a56pla4/7WVqf/tUpSfieCfKLZkkPWv056M2yPwO8EazA+RyyJSBIRwHp0
8BTnsBU7oN6eCvnBNAaFbxFqnqEyzds1KiCzAJq+/n9jWPuGMDZjcrdkwX1H6RSyYY6cl8hGxuiV
ZnJAxCeCGjEnKk8yqoE4Y3equQo/0GmcHKJdlsulXf2xucpEOcpmx3RdwmZONrqag3vYXsgGziG4
cTkDZkHZrdezFcBWLhRghgJVCjIPm/WpxIM7ih6JXYMsjbuP5LTVHHRRgmRvGyjyqZXIiaoQyDJ1
hC332MU1wODHX+xSYDLs44x5r7gMMG/LYu7FUSXWrLbmYGRB+3GoFjT2QeaMrX3YneIykb+a/FoE
sxRXrnBjxOqIlrPUCXB3YRwnAuI6q9lpXoN8smYUB0bNxwLgk5OjvtVzSm6K71y1rv0/ms3x0fWC
fBHzKX1idkK9eLXNz1b/Ja3YKaXf2qXtSuTI0uovlqT1sRM3LGbttCGh72PjBRpp15anI75v+5qs
hfT2WJb0V+AdylV0WBe94yQuTYx2+jaKaYJ4Vzc16A7tkUpL8ekA35uxTVZbcYHr84Nm06GwJ9GF
JszVusGscF+AD71FznEo/1BRIhI7xr9NFOIPVlR55foPH4jCl8tszEkdF59UGcSPXskOOMhpOpxw
kU1hPp3ZdJ7QBi5zPGtZYJdMHmqKAWQ/0Ebf4+r67R6jlTcbDkNYwXtsPrxGyihF2hiiEXnHJVxv
w9tFFMHclUKEcOHqvJe3C//H7c/R0/3JWI39DKJ0yMd4VanWgEM1ocAwPMMojLkVUNeV8hihOCie
/QYW2jph6CupWa5q5g/E+Iuyw4hfoHDQCvlYcjgu/v9uL6JCK2Uj2sdKYHrrPPJ7yrohE1uVVseS
o9TeazT7kUQDYZkmrySPiRK0Ibb+iqtGMt+Z2U5APXrPHRIhUzSgYhk76fc8KNLx3MG9hrzsFcvI
gVq00xH4Z8V/2MVLnhIjT0GBP9DODPgiDHoNO41vSkbZsPSDxMaIRxPQC6Y/mpJOdTlngEcO6X4O
59qtdqU8KTvJu+dImSrsSwLv3VDQlqT6oSXr06U4/ABom4UjkjSnERoLUmLRw180vz4rKaA1ZvdO
PcvVmfJzgS2/7oqlJmYrf4deJfHFFY7KsaPiS8ocYPVmQ+o/Pe9j9/nhhId24Jq5H/fhJucXCxQQ
QvBA2kHwdLVquxZ6M9zlAki/kWkXplzrjdrumzdWgfz8hi259gnTExvxWuh+YlkfP+EQYBTOQqGM
OqNKMQV7YzveBNHYbMP2B5spJ+C6fjxnS1i66nUdjlSNIqvOB+s4Dd7tErZC7BtlERWf73bgaL2R
AEUxuG8cEuToXtgMCr2TRoxbSXylGDEFM9P3QOrr3owLsOjEg3LYVMoS0WR2FImLDaVEQhd08ugk
msP8YQWxZqUNVqIensxS8VpJCn/nrD4Z+vh6HxP1Ki62hP2HnwJDiAVM8w2dNIZ2KE4hQQs6OFF9
1bEtewg0EstyfgUpagCbWdFWi9EzmVUq/hKVlwB0QfG/CzGRTBkZ8ZnzLqHpj+1EkmGQNK9G26to
+0z86puOZIknjWa59nWl0KykjIXUBvtuvJHhaFRGgynzUb+62FPzLmO8CgZ0Y9kgC/h1rbpb0oGL
ng5ymE7hJ+EZVRCmUiEfNFIf5k4kdXvgmenTaf/e+7Ww9XM86/NZDkQYtoJsRRKOUnYMgFREvHqA
Mn7G+3pKnIpgwd0fKdIYSLfKhQRjiZP3348VR78+pz0cthZFlLxBfP5snPFk5PrMYEJwrtcx+Qyh
z8i6WL48qJC0G96h5/ObkvUf/+z0d3m6x4WS6vBjsgfK1y6gZVv/3XCEhgzKEGX9aLqRiQMKYXhH
HiP2rCIGb+Dq3fVhNBV2QU/L4KAwnTJRR/Pksh9LZlpBshsJSanY1qvV7zV2Pyp/NMK0bz6Ptyg/
8Wg2cuWWVpiR3uyIbAKlyP3de4Q9EafTz5P1ZMYgNNo6J4ySe5C3ppL/rBXnAoonGvUpoAmUduHt
0+49h0yoV3J05Dwub+Rm1XOfIZzLj3QTYY8SI8gvXzJBl57HsKoD9r3Yd6W67/iRB4lfsZpOPPex
S2T9elSgUTGlIw4n0zWkoaVOHnIqD5qSCr0bvsLwhxTLvs23zCncnKH5cCYQD4o7vseRdxz8w+jQ
Czd288XuEV6e/l/4Wplslc3DXbaawa+Mw1rMLcKtqZOo4s4ZW26B6f3dIFOLpDG8Ts7ZrWp0JH6s
fOwqUKfFYP0w6eAjHLty3TGE7Gva5SQKRv8apcF/xo5K2C0VNZaqz7K6nT4DQKF2qYOJNDkZaLqG
2bNj9MXesaZq30MtCysxvcq3oLJ4313bxWwYSrQ25V8J38mD5y2idBXfw2eZcUqXCC8ilcbk0fuw
siNIT93ewem+ZQrO1ccVZMe6Vat8iFHzafLpsiJOMrptH10rnERzt0EwQsV7IRcY0g4EOZiUjOsT
yCmxIGmfgFYRGEyiuTfsGdU+5Q9Nq8iGWL2u9Q9Rivjr2bNVQp2P6nU5C92zIYlC58ojAnGiTkiX
PoeMu0fJLqq/owIoiSRvavqNiAVoZs5xAFME1HV2S6qLpBgvJwBsx6wLJ1PI+ZuJH3bo+78ewWu1
B00A9IDNHP/2iWGYKgCxPb4xoNLY8T7pzOJWB1PQwQHWCLvM9JJPHKM8xiXF+NWiJPkAyBph/1rX
HYtaDzDe63qE5fQxTrn8t6shmErrIPALiFZbLcqkXAVRqBrNMOvm72WE8puL+mKHK0Akr8cIVa/0
EGiSVtyTB6/Vg26AQqspUOrm0ruoDrmAmMVGjhwDoF+KSUwyqyyByFRD4CKzdtq0aXI9+85JjQGL
FLI1qHn69ET6js/VXIOVvCDLd4YgIkf2FHh14i0uO3pWod6SXtzGYuQqqgtIboLjJYX0HlbOzObN
ld5rB/XSXS613a/yJE9N9uQZLKQk5bKvw72uitAyO0ZcY6kKS8Rj+h7jWuBekptroKxvD8RBLFhC
5XJCXnM0R6h00WGFNivSKT767FcuZr/ZkTyM/yBGBH5vKpC9fJ/jjjN2gBdseq2TfejHx/XR3MI9
nqlUnQYLc5uxwnUjG52cB+laEQUQ6AosJKp4REx5SkWzKL6LHyWsoaSF8/kezpS/omtazZ+z6Eai
D8KdgwENHgNr5bae6gTmNc0Jwe7fOD/M7yKLSsZxk5AP1DuZ0/sX/hx7GTVukYzlmieL0KjwuRFb
PI0xAELyAa9+qiJZg03QiaqyNfSjiG572yPnbGShfOZJAwWBxstnYgyMR8omXrfKumg3MjBZDSyS
u72C6XqR6TprKpGwoscH5Cwm1qv+CY6q2Ai/ma7iH0hAz4bj9wvHUL39B5m3Pf8+KfY7ZY/kvOea
a/pnGCnyKlRiEzPEipJvU47gaAqV9RjmO5kkXvcmEA2eLl7M3XAXc4k+NaO7V9UT9soKOaeKTCk/
z1bVsl2B8skwi7iCYYzS0uh85q4J2mjDhuCVhk86mLS5go52fm7AJnvTlsLDEZ3gZHi6TQTJRDQk
6jZoCxwGdjnpJe7skxgsTZS+qNKPZXmeSO3XMkJVMf7mobVj4wg2/WkXHccSNiyWUiBf57t51QD7
/nx6eOAxl/VjiOfPY0QrWOmWotgxe2LpJVrKzQBZ5SimLtCY6JmOLU9QVagXRn8pmfoOwoZg2pEQ
cXhzgDruUL9WiCEo0hj/pzikzbSpW4hLlULah+CAhdaoW4DMvGdGY1TJQgee8+pRIXw0tZquV6SP
ZokDJ8oeLDa7aiazQ/OxOHuAfvYxKlVvHuiquM0zrnqwR2olm6yeaSFe7n5AQ1rRri+ReP/Ymp23
ympJnVQMo6L7TnZNZ54gGuXw3PHiKJ9G498y7Q9TRKpSfWIDT5bZoMphPs+iAhkYwe5MH2wwVvb0
oklpXuYQOX/kPtnmzIkv3G83lCJ9BK4jFri7Jow/sJxh7cgiYQKu5/Q2qaJHkYxeyUJmpqzYqnKl
So87mJGvcJEVmnvAyXUZRsmKKCokWIQxr30C8UwfWlquCJ2gLr8kY6cGEiGOvCj9Nu8iG8hcinoA
GUOCf5dJWWAQjFvJ5zkTfDkjv935Ciw0hpudZsqWLRAt9p7QK7EJJC3Gg5BtMGCbZysGSCYVxTE/
WUQFoWNE7GtLMS7m13aQkkK+rkFY9bzMr7/0urxSDjP36uSnmZK8mDGA1JKkiSWz9iPsu5/K/mLP
d34RTYdpS5PXVsZt2j1htZaxereGrnpBEglrACaZrWRheW2wQ6C1b2pbjCCmBSTrCS+temvbqXCk
Or44VwEcJji+QOkwwDhp8RPPNsS4k4V+exOuaYDWtymCOKKJbSTHLxC6l/2Fm4p3luBZE5SMkE6J
f35sxsGxDsFf1old5Fdt8CVXIAaAt+SXx9p342uOVtf3x5vDoCevFDkx3S4D5cjGpLiYCUYPdZCp
7dBu3RWhrIUK1xhuELvXINM1hfLToLQNwNMbU1uCeT5vRToGat/0yiNOHbC0DQuXuB4euyx3uZep
353Df0/aHGip30id7l9Zv0lJ9IqTZTUzdBxy0NNgRjCnEuQ4Fdml7B+A/E+85QmOF7xeGpB7tqS4
rFVvGazLFcI7ssTwt9DlaD/ySHsDr8xLnP2qpmuDSnnU2AaHFXgYj7gxjPQy4WU/y6yMPYFhoKdC
cmkoVr/GQ9r9eiC8ONdOhVmgkiHTslP5kyUYRS8v8gvhpZQglVK62dleXkvpFiISsuiDPX239uw5
zXom12uM5IrIKXPw3nQHdiBx1/5nU4Vi6MOSp4yGTSSeH+GXgxl+ffhpQ54kSttaCqCPpE4aC5Nl
KKRgnaRn62u5qeFmW+pdfFsvwhxKk1mMG46Xxhe1zaGQ5QSfTiUQY8QouMYd6Y/TwHBhrh1B/Yxg
QXwcMYqV6oQK4AXqA+GnMZDlQCBIt4O37lI+uKISF2WOEQldtu9Nwt4c5cq5HHEKoDWqJ0kJhG2z
6M6L8nGSsFxhKCtIVSpchZbRiDgsrbrA73YomFnTaGIbIiQSrH5BbyQ3KphKF2YBlNbZbEj5RBh5
DVwpFhijx4y28b5A9sYRC/Mg7YetLPxRSJ/taFVCPDQTo49VW9A/S21YWL9NNWuhMmoeZ1N5a5jL
sTUyv0L313xuohSbv2i7TWuhmmgp1vJwnJQPXwE9o8Uqo70akPR4TPLEvf/gvLTvfHrXEXUaxIPY
qEHjSufZDBfgNhYiYV5/7QD+h5uH4rOf7WM6gKgBlrU/2lrBgmU50IiZ1kRDBMgG++Ky0jQ4UT1/
EHm0qvi+JWFEoVcgPOckyEfZdT0PGlNI5+tDJnunJ2mQzi2TDomkUKSJ0Ioq3lzH0tWJYhOn/1U2
ma2HuQB7mWXHfj+/ndmMW0nkftZjBd/yUKb4Pl7TS/qQJE4vJhBMhXFMtGPRv1svkurSPu4QUg5p
owgpXjdw+MgJcFiWIS24N5sd15R4uwwoocGeIqYhCv4TPMvlt/zQMdK3zPXxfH6YGf7jq/TrrpEl
PusRBN4gkw6K1UAkMp661NEHhOxKgVt0azWXbJy2wxaXZMWc50oXw1yhhil9ishwWQakcee4+xr0
wKse9Qx2TR6hWKaXOqgxxsSeGWRSm1XTC3m8Pne5LTeIOuNQ8AvAe0gdvjVManVV8EsrSugH774j
HcsadHKJ+z1UKxOAfjZT1qK7bJz4qZhraZGXW1cCcQCmM0l++88VaNJIeLUQJJ8KwqxmZekv1USI
NKeJAvR37cSXWxIr6/t1BeeqkOr9C0cPZVd9GWVjpqdggplsf9sw9UE6n1IvrXHZFfvNUZtaLt4K
W3UgC8PChRo7ljo4XJL7k9VFpChCLyyI3S+X+hkEXjFdcN6obqyskHWlo08H+XjkLrR1vM0apDep
ggQPro1n140ktM6CAx8N4JICEcWP8ZOVqXqrgocawIzM/h6RMGSVZTpc9Z5VO9kGSU7U1cbp5plj
48YjmGvfPc3qYjV13l62YhoRd+KJiMXs/6fUR6EsoMM6/SyOKM7419dlMxB4oDxphE8l1/9WEWq7
v4oUZ279VyYEMvMI9EK4TYadWA1upIsbM3em9auG/Z6OHXqcsoP0svzdKEQeA/VLtdQHz9LVcF8U
EaRUlkeET1AU9FoXNrLKkPuautCs7E45TpfaaJPXCeqgOlw7kXhSdlfltePWwPOI4SgCJhLV1Qt4
REkIVBH0S5MjS8k9b/efTNHQBuaE1k06qODbx2GcITMN6nW6LwuSzMvIpY7QeoKbg/Ckp/1pO8Dt
jYub1f7LOSyehZQWMnXa2SUjuBWk2KwM2vTnTRb4sv7l5vodHeMfipJPZt9BE2dN86AJtOLAImU7
Fqe2xCX7se6sLmULBjwmTQGLwtznoWvVdGSqMz7Vr8A1RRT2ZJamc9DFuckoZ7J21I5fTyRN/mOp
ZFoeS6yzI7/SXoN8QjI7VGB/9XrgrwruSeFnCDOBEpaK4e4mzSXWNVki047JSB2hvILYK0kh79wB
91ATo1l8yuUUWU4IYK2cOlA3NFmyfYxEOzlnv5V/rIlxHHu9hEHJBsi7FSoOWQdhkGLEDP/KSO5L
z4xEhsf0vG921VqlpnA6j7wFuPNlqzF4taJUELUuhQ7CtLOBdO+dOowtVbX068csOGLxgEfmvtSI
fLPDrETkUkWt8M/yoiOxDt0iJdI/cG2fZ9dpuBKk1fsnztyqOkFrG94AZeDFyXJBrCcVAcrL+f6l
Xm0RLnZXO3Y5P1ZjBywdiP9I5iqzVqoeEgnVTV52bU51Aa+AjnQdgCErTFBGFzG1+HaYuzNIdkij
RwbDUWUCBCEZXO/z3JGXTmMhqlLF+7b3y6M9vNZJxEvspYIJcQj+AFUwb3mtcbuuipv6PIwW8Zqv
clBQms0lWbDjHQEXCEtP0ToetN5V2owA48A5jOYtWBVZLEk696V3E8UThf43jiHpLb17+WyNVW2M
FE32Ct1Ch5WrdKyDj29wFUB8qSwfLdEFxyXvjPl2vAMHJjnYYZ74UWm1+Lfv2tuO6ZNU7VzRpZNe
GEtz/m/Vd6fPlktKMs+QGi6NhAfeDTRxJojLPaQoSvHoar7AFwmo9ODZcQX4B24h4GN72TPmFmw9
e7i/cHKv8ie8EVn535cw1YlcjrR/AJVuJdO3XTy6XqsvHAArrly6mnnVgIdsHfaOtaX8nNLH+zS8
oUF0UE2dg2uo4ygx0wNOiPjVvrc2d5Wp25g/FJLNCQy56wyU7cXvg4+UDm0/Lp3Du597TJGSTlog
TQZTqnbrSMcuNFEChRC1Y97iLyFTZ5giI0BljhIDLstDifIHaRvPb7m3laqxIQh2mf8s31HU2Quf
I0PLsZMYFG4v/01BLYAfVcD7mt25KRfdlUBv2qMfAW1QmqpF04iKLQy7sRHlKaLBVTeSfNHwxQJO
sflgLsUB+190KaZ48/T19WPPSCMDc9o4H7ReLPPiLsvcMLleQ2UWL6KDhr35gEdKhUQOcYEgxHmW
9P2ll+1eChVPKpl0DJYbnjFQl7ai4QnKgt/XYCE24dFhyD36aQDJ+STOGPUfiwSyouD+9YvuyPX1
VRxxW7YmThGgBcFRpechti/8J5FRYW4FTtO5VEwJ4yr8ALfTW6HGJ0aF24YIRK9RbK/IDbgOS300
eARRgSTrPM+KlaoUPbSQ7/MLW0KaSR8s3v271Mvh507LhwMxL/EcGePNHP+iRc2/P6r7sEWoeedr
7GPhtKgC3AhZ7NCg4oCIGPeyxRDrAYobdPvpZYjP2jUpgPT/E1xr9taFiyjglBR6bKrNSiaT0b4s
+7litt1Qz41QrC1CJU8iJEMtZkAk4gxNVH8oC/CZi5jXFt66ooixRdraBkbIe+HYJqL40+ISbbgg
aEmw7HVgA7orViEZ8MSh3pdToCYQWIj7Zh7KMaILGWq2EgkTikWnSynYO787TO258oAel281zbYA
nFA1VNb95FMXh0CqLuJ5vs6kDIenbl4gc1fjqzKGw/XX/BWMQsQKS9bCIjElvi/dujfnngVZIfDI
eR3p5Jtrlrs6Z30PTs0z4xUnGQmmXMpkPptzIjoHYjukPHA2bS+oNlYa0voSQU1ARHpC1z8eokZq
zUWcqp9IaXy8uDMF/13ZjNUzMcACm9Y0Qo5HcRv9wTyf81ezgaH8pqVdeVXKkbSawCqlVbCwy0DU
+WqCYkYSeDDlF7VhvqNTcqoCqdwC3HCafMuNXByQ5VfwjYNaWU/ME4EmBBB6pqi1DbkQA8b4EOvR
MsayVMugUcbrv/QDg27zAU6L9q9JaOoHBdaoJvMtBq1mBUKKaWJFfEmXNobqL8UKmKhgvtDw0bLW
wCdP/eTqIXoNMatVpZyOX5xg0FJNdEvMpW2YbizLNefECp54RoCXESLg98tWX3k0ZkkB5WIr5ZJb
0AMf6m5zztAvI3sRssCH6bicXC+hp2WP7YRsRyt3YS2hd+OjaogOFbW6WbBbUUr2LuBi5x+hBUd7
+PtKdyIogQl3a7MOaqpOl6lvpBM5I1iGmmYFo22CO+3+FoYXZLQmqb51Pgc3LiVDQcpJpCBZRpj6
KNjkMfGzUf5ATIx1HIGFEiFD646SC1fT+QVc6u+l/rgeh/6p8WxnLblok1sMpstS20Lgg7V4JQ39
KKx+6jLbksbeZHpbPRWs24+yGmTrm3IGvVjI5NH6Mv1t/Ez+p4T6j3eqbteVVmR8Vm8iRe0F57nS
pevO0JRlQljn/fDNkxkCDlgODVwjn4fw2dt5UxJLZUMQbl4Cn5Vo2q2kRBIa0LqgzyBAujQCQVE9
hRHYVKm1NN0sVYhGnW6iXgxUIybtgPqqwvSkVX7/9VijwzrauQPHx+dtrFfeV2uba88M/aMmYgrk
67RgnkA3mmNfHfWcMUpWahqLWD7dbfgJO1+9d4fubGJsnjiHnpxv3KDlj/TscHEO2AYMBQ0sCmh4
nWFOQ0v5vintT1DM80BzL58HkOha5VwyFE5jgjBwd6H/qatgoK059qVg9+gaxAb3KeMuBQFMGh7W
0CktalfOu+jbIWDL2CzIlUEm+Y77hIpZZHl7cu/nnl2A5ECBRz6zeTJOtZHqcMgCcL0OroFfr92O
EC8795bOcwJwtQlriiZZ+HbHfoWK+8Ao9w5Vb2u/2bVkhqQWDsbAtCiUAi1NtrAFWbWYMBefRfCJ
6PtYGBAKAASbK0InIycw0bxdY/tcZc4hrpjqbizoZlKKX/Fe/xZdOUsj2+4jQDYobg59nkxKczij
BU+0xqTcQipwBcocM7/jvMcQtdi4fMeGZ/4ZLdUWUTB31VZ+lTFJJruF2v5+ML5Pkv45I/9mlDc5
dr+ka8oPne3GTL00uVZ+cMuYyoAZnDWdPXGjUPeCotYTNVret1Z8bXfv0THnzLGf3K+Bh/eRbnka
0TNyltCArSxUX+CZDyibLjpjZOoUhc1HZtUcqeTTJTSO6UpI/szeRO8+C+9nCgyoLZ0b8puhY23p
0cPxSTYDKumw0hlMJIrzegGQPVisXtSwDLvB31gx0o1OPsVjisRK0GGDXB5NkYJEGvemksFTd0Mu
Scn5j8nB50HSuAMLJtuLkXH7TVw+vG9UVroIF9qOXjxRZVqXxcNssbmnSwwKGvaGBbqfyIfImYim
wROUaREGOyJ3EAbZTGdlxQb1W6jAOMQAvxvC6jGNbFulZK8xEbUngq2JNifzOu6meUUeq0FkT/am
WCsGu5BUHPG7C9awL1UVTymtX/PZYKQrSTXJ9jwegX1iUfISERXtKjV8tWb96u5VSWMW4g576PHe
UAEIaTMS5QsY1xl6dQdutvFdbTFX1gbEKmU1ds+q6aiUUZ+lGUXAyoOSS4AjYzkgd/kKxyzmEFiE
tTWcGmM/EdPztNgoHOGlZNN5kbVLy670JrbKbMYg9Dje4RdIVH8QQMkyPncDaTF4sNY2yBQQTWiY
HhM9OAHmbJmSrXcNTK91kihFCUlbF1zUMlUzFdLPKcWi4KJ7LLQfEEgME6flojzNQ/86reXnKvEu
S9RHozKgSbUIrVdjR4Idm6e/TiuiWvZdpBekmrWSkJo0tnK8QSVJT1BY/LR4lhLAvY/y9OR5gZs3
O5CXRER2m7ZIp5jK4saBezp6/ekaZfjJ07g32+pkeNoIZyLO5Rl7Lw6/ZVkfdQ9VPshyPhzjpMIy
xdaf7mC3SPZ2cjpMFxm0HphlfZk0a357Udt7LfOfl9Q5Wh3YvPpN88Eq3bURDJSeeFxfRzCT2tIP
NX4Pt8+0qKve1qKkjwleh/yZYrEurBJsrJyefedOFeG5s/zr9eYCc0oi35IZuXfx4ZZKoWr1H9ER
S8/VtTgTAEJIeXQRN94dt0W6z/PVmW9OoZNXtUyt8S7dqACks4VVqVIgp5qR62Kxb6tpkmn973WP
Xq/c/IgzN3MRiWoE4W3kbP7psZ7alB9kKvzRyI43LPzeC2l8EHDcturEtp3ecV0/khkMYsRI/UUy
wBaOc4xvZzBmXWzM2Olu3/1ZSSqA0DNKzAhnf2BurfO4KJmJZ5d8/Fzb5t/KBz6UfVJaIpRUJ1bV
q8iR8QHN6WXXfZvWVxjmFJvsP6/hORyL/BC4jxf+Yd+czQW6BxLEfev1F+PMBp93yHSta64cqQ/4
Ula1vBwwFNWvtO0m7objBFocv9MvER/l1WZa2jp02afR8akbugaXr9I666arvgY1tu8ZRz8vr7M5
GKtluaLH76pF0KbxBE5/nXRN88r3HPnDZliMjvC31Gc8T5ILGSMaCr9smevG1x64Wk+wJ7qeKGJe
wPsNbft3fQ/wZwhzt03b9EJBIrPbhu29ItQo3gsIbIvoj9GU7ncvMmJEfrSI6LjSVhLw4vOc3SCA
TgfD0nFeASow0i18hDwWHfufRsGYbI9eHdiBe/4lJKMGQO0uDmgTSwG6beJS/VEDjxu7+Xslfels
xP/5B5AdXjtD6RkhSnrCT5uYofDtmqN5CzrhIJYk/sl9V66dmioyJQjjdVHG8Qv5miUT3k/7+2Tl
BJwmBrRZ9wc9fE+f+PsLqtRaYPiPVBuy60x+pN1YacyroqA5Yh4Syw9lkH5tyKimQCLjW5hDnRpj
cipZxuy2GzttgOVIgrp9YMFWHR72R01tYHQoe3AucjUrntvuRez0pMIO7Jmq8G1JFkqC4c94axR5
iBivOVyry/RIYMOnONim8CG+IWhRswD5m0RSqj44/HSUs9FCeJ4HLz64ZN5bLOqTID4yvpXahvuB
6llJ7g1PLC79K+ykpVW00v1O6n7onXzxmr+vqpRYeUqpgPQS2HZXfgO3VTTHULAI2GFfGhYwry9g
8RmGhkIiXLCzgMXOCaopQMik6u5/tKRTHKHXBcCkd7LLr7g2o2lRyywoyOKMkbKlzZSHuYwqLi7t
yuHs+JivwlgOAc0ga0wbI3BApPoU9tAcm3WkKbSj+t8FrMaBTKA7E7vs4Kg3N0Cky/lLsmnMZWwz
jAYs2pOVNWYv1W9jycnzuz6FRGBZzPy51tD0oAQEIGWzVy1wmHJ2JRFodJ2Lc2pmYNUFem/MrhTL
c4X2G9vXDi9rAFKAMIyp7ZWZYQAw6iqTaloffWL2Tl4cqjZsM/c9oaLwkkxtrv4TOdglI9A5N4vF
PKO5T02gqld2CrELtS5m9q0Hq3E08M1+1xUkXsrZpzLFuUyWBrJP1QK8Y3LDpxcdhpy1xk7EMoHN
dCrGU5EoRvmJYWNR/ZTDrmNyLcmY2atRmUQ7+lX+RX4kdnwuo5bs1ktXLpg2DZc6yKMVhi413ERb
mTYTBiZ9aH6z9CletPmOvQ0Vi00pCFMEToAs3GAzQ5yRfXFhOw8aokz1kYKxuvYu4a9+ACDS3hBz
6BhTp9LptpaHTwg6uI6MD5VWkv6w9PkbS2RMP57+97pyJMQLpKkjsse6YiaLB2y+IOVhUvYiU0ww
mN06JUwJHJ8C8z9tImT+yEv2rldQJtFXxKg3B6RmcBkEz08SX+mRda08XVp4ZOBIoGhTzMp3s1nI
ZcJowvQtpgLeDuJOjcXnxBuPYX3hNiWc4ujsBKPuRppWhNbEpHQ1IV+6jAYvKBdCA8kgVJLWwJTU
KByfGqxI7XDXs5N2uGHbRYLJ9NJJ8b6/YTM+PlDgGAIbJc0DFLi8lskjcoD4k6AMsBf74ZSx6tSD
R1qSeChMwzuVN8/DDDaaPC2qU7rEdf3xL+AOrgHoDW+AUUV7QcWRsZaDt4laj34vrBKC4dEa8qz0
twYSA+/L6hsMQ0kDd/56N/8TLJvTR+3zG8MJDymkgnOEz8A3s4SR3wjO0ZezSQE8UbbxMyewQcXo
mEwjReHaOImw02ZbbGLU7TbiFV2uEmRC4Rr/qb9oO9ZreZ+7sH98O4pdnD7PfZSkLDKZS+L7yt8N
6Rg3yDm3EPSG/TsKMpO6mR8vRmfNKBSktqx2Lji8m75eVFvWv17Zbqcysc7lHDUXLhgT5SU6WAwF
hXhy08uuBpcNAxmTuKWMiSzHEJJhVZt6oA2OCicNdwuVpdHlNCrVarujBNXAUvRXGFpJP9uGqNqE
XuVdeIYLxucsLegSyAcA6ZOzOcpuaAvDQp/Rr4YAVxpgW/Tx/fL+EvVNlUIBGPuZm1pa3YttqHKA
CINbvWgk2HtwKcxbGQuNFjkAKaAltQCTeb9yT3NoqhG3IitpomQf7pebTKuEjZnAJ4o78tx7WuiR
erJryxjbZwmf8LzJIcpeTV5I6L/cn9E4KIaVYfRw2IE5gHeoB/v+rugXbeaqPySMwB97M5O/Vjjg
fmuqJ1M4K9MhEs76/F6KKBTd6GSs4pEtUmZVvLuuTbXECy/PX1wEnpifFHFGngnRKHTEujG/tz+a
Q9scbxMfs3svirw1Oo3lnx+7kpn0bDjn4xn123IAPh4GFLdRvSlbV7fCF3NsVLepQoqFOxHs2KHl
I4Hz76MGIUzpR3Y6TFuEKG+CTgHcJ58Mn8YFj5YrVmUPpfFnpkXc0o7DheARzetK4TtgVmFltDsk
FHZWeyU0rZ25JgfGCdtTLjqJT5YEjrbqXmaXbkKw+yHVcSQjEQmEap1npPRcAItf47wuovdfZNPh
+RwCbj2Jk+xC0P5MTktI4SpAseeT84TPDG+BPX/zE2R9tl/XQd/omvW7MC9pulHtdtD0aXU4GrsB
y8sTGAUyUWMsgvYnDi6IYnZ4WzcAF7cByguDolztn7DQKiXyi8NSnvyTv55SsWGfPkoiregk0LnS
ZZKtyQs6rMizKdCD245c/MHZ8EYW1oEyHEQLPCvi57PVtmmmni7jysmvSBpZaFaMqibi9AEVTPiV
tJN1QMsLunNQ/jvAtaYz2YQ/U4QPfxXhrjpwXYoMsuBil/Za0/j39eaq41WczFeeMHKAJ2kdT9xH
M/PfsXXY/4gMJ4LaDc5yWrRutuWJcI/qUSLoLl8Du8EMUgmGknfNPw/F/tblxjbQ9j0jJrV59BAf
dSI9AxtjR9b+Q/GQFqOQ9WidLTWO6QWtECul1Jf1nK2oUTXtC0IBaR9q18AjxY+/iRqhESb4hYVz
obG5zeWMRYcjqpZaEe/ogudYga5LLdARThRiuvlM2pdWrax9Nc6jK6HhTUdJ5jbdWm+Jy26fIqHO
mdEmbS0Q2cpaKyRJsG/8NgwAhFuE/JJLw7ck8HjEgq78YpL6QleZIGrzmptBVvqd5E7NR2mGmFv2
uIE1hI0eyQ6yKRmIBQbS3DeA9WojRO1uYZi/psncHqQ8IllBlNQMznIWWc3GiZhzP9KhoDFKRL9C
Mhl7tAOAiUnI/8ieLsFDe7Bd9nMTKl/N2hAv8JoQ5fvfLW2Gea6yuGp9RuxT+2+tOEMhXEgWcNbb
PR/C161KDiGyJsBvMQUvZW8xeUOGoALsKXjW/jrwxZOnpOc9X14JbnfyGigiMsjKw02fqMBi7vi1
qO/qHIL1YJxiFWT1BWDQLZwzhjKC6HcvjnGxTuUMYQT5MpFIbUujog8ZN26CFyjeOifWpqGy3jNj
11FRskDxZo8v0xxOR3P8KPppxTAfq76jmc1UYrO6jo8Zx1Ss4rsxMb8qYhaAHCwYZAmpedI92oTQ
t4fyKZ9z/kmpjr3IvN2c583DLhZXacDV0UJlwih/MJAx2WRJkmTFjO4zjfxCTu2tb4lVghG8ZhTY
cZmiwRuHk/HcXpCMAsGcF4qpQEbIfNCspG56cgbAmOVYESc4mBI1b1L7nYg6mYKle0579Inq62al
NAaKlsmQMlBoInAWReptPtSNKSt+m7byhh5C5heSPvwPdvprNzcFzdlwZlO25EUbZ26BC8/JfA1b
03SxN4dSYOFVGsXdFLUqX1WtJTO35WXD9YnSJ9j/o5AOVmkbn5JzkfYmTclbKqcLFD4BQcoKDOM3
cFWmeJ6EbWQhHqaEsTi4CJ0nElfmsfpe5/dG3EbBd4LTSn+nlnRuy68uy30A0n8vmHzuLyAE3Oi8
FY40EAQvP4nmqs7svPvzaLrL1L8CAuyVTGHk2HuI6GfxjDxQcf08J29iAPHhO3oy8QG6/vgf0AvG
TGrlPp+AvO85/Z5JzGCMiVKLgvdQoAIDjchnZQvOwWA/SBkLEClcbGgQO/3Qfkq/2yebno0UBVf2
+S8KNIjY4yGK3SEmurF8djIfDxydBu+LEJ7EFFi2+YM1/nAlc04xbTSAUm9+5tkMud00gGmFpA05
S730c01xutdGBUW8IDyoEyaasbSTkJKqHZRwC+sdd4prr0ei/xbqptrJy49BCkG9NAXwSbi5jghh
df5N88N1ArX/AZHQiJ8ruQRbiwAEohHS1IQH3SftJCk+LXZ0BERgaTBfhEyh8UOESLyoYWhmSDfR
oU8R+MW11FIk8b6DMH10OoZ3mQy14fawQ62FvwMVXKZRQuk4Sd8I7OxihvFuR+Jou9yswJbXzk+o
S0ZyNLVxDTKG9DoN7PY7i439488/qpW8Aru0sJHxhqOLi4qnhBoJnT7haGS5jD8/DSvATOk9f/HR
Gcts74d9/TqblAo+JrF1BYX4S7WPGbL5dlfAiMLOu93fIauW6e0JcLSCpNx/+MNg34xakAqrevJ6
AM7OIdjXz8sxM3ODgkdNYLiFtWU9kvNbC/sE4d2/O96Cva+7PGcxLaCfSGCaHzlgRn988SLIfHv0
/xGCav+eMmF2YyMtDkikfpY4zZjvKnRpfKw0VtnrZ8w/9L2jPMsE87QtJY1AdWBfZbi8l4sdV3iP
Pf2e/xX6aX/+KmFuDpwB7aeobesDVwdA652/gzusiL/hz2tOCb4mCSTeRUN9v/ujhhwGmKHoi+W+
LODyxkoHtiAqbNTCO/wYoRJ29ji3FNo3OCKV7eB3rtZ4ALv/lcs3Au/EI/FAC3v1LABtoUkzwWu2
tI5Zn70FxOq622GBcHw5xc4uWC+oi2jtwY/WW1BljnOgOaPkqU0GLmVlE1zj+yVVcl7o0eOUngHa
dEB+VexGTF3GEL/lIAUc5StR0v9o4VMAWP2eAZ8OouGPysESHncABFoATM7adxJHHRwBfwCb2Zks
xvqQs+gmNLw//pibrZOfsVRKYXPGECLsInLazd9oEjkFhVGa4e3GI0G7ZIQKxJmPuoTao99Kh7Ia
ofvff6orF5pHjxf/mx/NolYvsmZwTuJOfGZXifIJ2XjWtl5AHoLdB/IpsVlC0teRFw93Z9gfNtnK
/q5+mkymj1L8tUlrSeD3akjK9qWES/Y5UB5zlfSM18+koTz9z/it3qDQW23bzvs8CZ8ntWWOjdA/
qMglR4TFVypcYYrDX1OVN5JSsEoaUkymVNPRF4ypiJH9VFjcVIUZ8fB3iuz7B3DDhzpiadYJz9VT
LtuLfe10ha11RisTxJlg/5RPmm9KO0LBpKDHxmnbuO0GZrFh5mQycSK8Xr4/+GSYnJsbEcrcityW
YXgDixhtrzIIAzePR/kbFSkms0uCDuGoI/kqmo4AHovNbPKfHcz0ZSuNIy/9KMEiovFBEiQRmxdl
TsDtHP6mZRfIfAD3OI4c+lQb6nem7cHBayhA3WxDzZKdNzo8Qhfk/WqcFXqfwaHe4C8wrzGRCyM+
MYBNHxQ0H3V6WGbMFR+OWDOftQgxwoc1sH1xvE6uM13ZrSqDxaCF/WdV+wTzmaYH/2q5nvZkt4Rx
Wyv2keKNA5P4qwtLuKLQBde3daKZVNhSbgizZhblEbLoJk8RPKpsrt9m8JTlKioCk0AjFwQivp0p
+vom/YJDxLyKFKLStxUnTW/m01HaGqmzFeCyknWb5yN1Vd4ZST2IgsTuiy3Iqh2l6B1rBLCOfrFn
e/gDDse4pPg+jZEBUCVlIxJZIIxJkDZmL1omvGYoCIYjRwPJhlQfXlB/eFDHGrVqOC0iiT90N4rE
dx3prh7Ze6OfacV4xRAQG3RZvChP1T56r2gL7LrJa1jiy0DWY/9T0CEzibeR/yjkhkwTWfcUlNWy
CMjgT2zNawPrK4Lt+85y9d9dTB2H+ODTIYJQvu3pGXf2Ss7BAI7d/xdN2NhjE0L6h6GvX4d7xj22
3JuZmsWn/Lvj1Q/EihRHTOKQVUNMC7ss9JAowZsb6Uc0kMSyBniTsbP26EmalqWdu4gKOraXxfhF
vuvM3YA8QgksQKO9bXW9O3eOqxAtSYCAOu8ISf6NCCfN6Yi1RBUscHnnU5ZQWZRTFbH+aHL3HGGG
/3NVXI3KHouwTKrzlgOVX5PbsEBh7CkuAjO0x+nVH8jTP3Fjopm06ZaWU9Nrtg5BzYdAEBBEaD45
9KI7ulbS+BL7EhJHBxAMdBzEepWPU39RzvTh3n9nAYfIfn6wXGiK3kCHZ3gm0Wmzy50R2tw6orVg
vUR6/FxAkd1nYylKthxjCmmE+det6gOcGEmSzcfSVGTa6Yegx9S/hWD6IDzJSiO8b++9kA7t7rbY
zRqdi0mfzawYzZJNTjKsB4v76beNoJR724fBryPfzDXxQak/5GrmuqPIuB4+cA4F8CrIWnZdXSq9
TrSi5zdXktgpAV2uYgrnAhX58G0+8Ez9DBPY1lHEBEMO+1DfpeVFojWGpGphZiVVyELqt4ub/Jlm
sOjQtGFip8Qn2x4PrFo00cDMGJOkMle4quJKA0xnH8bJqpJh1xc3H21PfdRAK1tnp6PnVaVfFuCn
dlaQpK+/3Nyf8tSeHSDg8LCWKPQDJbpPKTmxUOFOJhtygXEM4Dfg953rsyc7JCg6QCrkPVmSFIIB
Z9fXnKjjrM0bcDLmOGgcsnQq7OEjmaqvPoOtKGH4ykTG99fWxrciQynpgnFhQrXojmJsre/S9C68
dJ/i4o+g75/YmLQVzNdSydDKFBjKnEzkI19z75jNqK91kRbfS/yR/bvip+qMRFBMLSrqx6p5y1qp
xmHbzLYqocsiOQcuVsnMezXNRMUWjWJq7HQkiyaJC1oXxt7rEXHHXnHyyY3AAH8UNA6exUSbRFGy
9PMS28mu0ANFe0L1xLEQx0l1ycBhQ2uDgcp3zZPr6uVUIlaXNVhX9Cd+mZG0Mj+65REfL8get7Kk
L7nwNZyZXUj6gjC12JIEKB+r9aUzwx2RAV+rufF71Ce+fVBQrq9LNiCnnTBy2eRShFa230MNAyDD
ME4KPIUv14Hbrb7vOkYWUzZQVpRrqmdUwqse1q3ZJzRxuL2d8xIUV7+/Sl8We7hIKx4Mr3lCeENe
r57azmIeH8t6zw6mid03W+mBr9u/ItGombmvyUh8BjDyTwwGOitRwmKQ3zBZpfbSIbwuQ567owUf
qRFEq8xr0VXpNAFC5ShV4YGnfi1GpiYMpU7DqflEJ0KmKSJywMpqINZG5IYeNh5V4sPYea2Fttzx
HvujAQ7l8dx5B4oCZE7vhtEhjy4M36Ga8blPbJQFHnV6VopdEqJ46h0fG1Xoo8cd2DtiwZrHTu0e
ABE0GKBCQoIgeEqH1CKqB2GL9Xp8GQj6J0DiCyuCifpsKELUIfTxQ908Wioc6ngwxRZoGjisKrJa
pK1rTQXOupCyjRVwPhLCeTwInRJjv1K27ApalY4Bto8iOmPUj59599VUgqT8b0/QP8Tkuri03Oph
sjT+ahkyNjaffwcKRt9boVE/1+FssD03hq3V6dUqngQK73Xqv9/t9xF3DxCxMmL5IESZRrfSCrv6
HxWiVq+Ro6y4BX7oaay3sQL4uEClKx/0FV7u5bbajCDdhnPIitpiUIpwTloymfGcJ/ElqPrzeeTw
LQc9Pfn3sb2B5ZCWU6JThbyq13SEpJ/KuTyjySJ4i4DIBY6x/mPaKy4bVKZeHOHUFBsc8L9Qo/AT
20/txA0n/4rEsb1R+n/cC1+lF66qT63IiiuzfNze6orkqNORp8EGpalhR6pfOV3FtVQ8pOa2KE9n
SD9Z32kixtkbENYQTMQTn0JlLKX1pNGRI2iZPIwD9LoJ1df+838qmWAbu/1hl5P0EMHqJ6OdFaA7
H0nZ3YcUnscfUzH5MFJQ8jo35+rGpPngerj+p9ebuqD8vh4dPTJMl8gntr40HcE5pbqDhWdwh4pb
nVKaGbyfXdFjHBlEl217qR8RCnhW3iEdvz63woOpkM9e0Y6LDfXQLNdQ0ENDxJouIJfWdmXz/7fG
wITB+Ewf4RFmcaEhEYd4O6s3PXqYxD1/EEvbS4f9Pv2lBzTCRDtpatQJ/FUsK3WQj7STLqrPucxI
FqrviU5+ftRfyAZW9u3ZcKRtpkheBMv0QamV7LfvykGZAjWSxBOLHyp0KB14IUeaUII47/souqQa
sKqckxXlfd6QchtDaXYFKJMVRJiz8WxByyFYtP7g9icLi5YTWz6nr/SrGSgKjg15e6uU2Ga0OBy9
EdKMUq/KoOX4LVfFBEwjqe/h4TwnQQ/Vx49xkYWyW/22e5rjXAqMxYqhLmY3AD5O5CiR/lSrVe/C
xSOiuOqfFz2/8eavISeinFrpl7otnawFstT2R9sygml4H8ewQO+qJr6UkwFWP87p9xs7oAdc5HgL
bf5M3FSohIfS2kj+G3uxOnb/Qo9wSEhD+oQ/cqktRF+ESK6i64ZBkGFaORP+u8I8244/UCX5qzfD
qXgkSZyLrdMnwO3q0fz5ALcoEEVAZ8XS9zWRSUSEyIaGfX6hXWJ68Zf3BMxWmqDb1I+m5BFCl8Dx
e4YDY7JHmca19SXCaNbt1GkrYF+IXFYUCW81kWYYxNmDjLM0rG9JzXBbLOnqp2s3/wT1P4kyjzDb
ZftPYc0V0gr0LgZvMYoH4UVN2hJWd2JmBlYURx+xHqE4l3jY0K6ylruMNaaNDDEX2PcdBfk/xGgu
9CBmm4zoGte5KmKp14V1IUhciA8858c8F4vlAn9daGUFHZ1cPzfKjnC+GQ3EDlJDaOki6ee5s/8k
zNJdlr+8XF+VIQ5cU1ZcIz8SQj4I6q2dZZu3LF9ZXls5oeCfFq59TkL8DXiJwEUeQ+fE4PSiijTq
rxWMJZd25K9Ww4/dtJdSDCMuNesZK9Dgx3t+mSgxtZo/Uedi2MDy8KGh9ZJTMXCoFhPoyst4Y/c5
Ao7Fq2GNY06YQ9fHG9Z5PDfSml3UI7RlRSHp8oGqaDbCAueStIgilabL2Cdjm8r01eqSLDpRHkTU
LM3/WzKtHMPCEpsNZIfzsf5en2+aViEw5lrlqB8AZsowquPRxdB4yBW9iG6J6SuODLzTi/h3CW6j
2ozSEXqep9ECPKZv+9OBfx8ITk+D0zkKGJwJtuN7Wdr0NXbqWQd2RD0ZCQ1OtsaeqgV68irKJl2g
ATa5p15/th36clpOnMZId1Hjyu7nRG3YlOFldsUgLSkTWV9+ORyu5X3s49JHUzp/15Ydj0MYk6/w
f8kR8M4gpBbOnTvFH7IheqkA33/cY1HiwI0ammQffH/NnYrgYU/HFG7ci5hx+xnR952VHL2fgtX1
MX8p5NNJcgvR03IoDVST+cyk+iykRaxdrDDWZNDhbfHHYkEMNgt3DD8Vo83JG3COB1uTBWDUur1L
nqQTW4bvKtbpTDGlZAt5j4ZdE8RHfFTbrv4waFpFqIpmoyDpg73FIqWfpNnBNtI1BwW9eY7oWqOb
586Ysg7Up5ZMvS8Ph/ymeDuETy8ambemPp0HuElW1zn4A+J7o3K0ssjpp1IkXHtCe7FF7SPq1VWx
B/+/7+oB3nZvyHAV9P8QKpiOKfS4f218hbpIslKDxhu0moGfm1QF+oRITvICbRaInd/0lP5Xefaf
zb4YuZ5C4h+ZopnTjvenXGADBAuTx97yqQ72N6gAyyjaf+rLsZk4ZDuGKFTVkeLoiOv73jgBys1o
JYuKv695qXbfNg7YOMgspBw67s9R3a7ENuBQUSXZia65NmjyHmpU8eQd1T88vpWyCNrDTrZjDkSa
OZmhRBHP9VbdZh4cWOz2OR2j1HXpQ9GAVRjS244AIKeOPcPdVnY1IVVC1ex0Sf9EnNNZw295yY8s
S30bwBUK46dcBuyIDYIGurkcBz7m9IjDtryu9T3Uan/qkf+aLCAyN5eaxnBRBkxKSFRKWcfa/Y+J
0OIjf/eA1fzNyztLVdWxEvT2B0fLoyiwVOBPtSPbVp2HO3qKKtmYrFC2jib+PrmFgX9cie1eEani
BVszQfpyFffxiChHpVBCAAMek1lf6MF7sEYr5mYcYoRmrR1j3y++7ULgjLwADb2+2Hm/M2qBGF4i
YirU19lJQVaFs17dmjm/h1hS8tlJM02QoVj6W4iE0qpc5HGP23LaIq7yFv5m+GsrFX6DfqufBcTl
fMsK+SCfFpA1mkauB9pEMBkRyUkNMgJccaC394vEbAx75/EPzd1fI60SeiQRErFFy8bB+j2lOaTh
DSQ4efyNVmVRF+FnQo4sMMU8AFgcQ5k13mWjELQhfI7PBrNBCa2xWvAhXdS1n/pjEPXK/16PQO6E
51Q5Cy7pRhZe5EqTjtTUHcKsdeBwZS/YNcDVxiv8mJAveJC0Zc+yCbUyYu7xqrI87q/NUeLN0tp0
aiXMuRmlwRIhaSP8eic0qUsbgDshUOcy4zCSMQGmQDqN8anhYAHoqewj2UeauRC7s/GABTehSCo6
hBa0rJDNeMFc0hzXNq0J6CobK8zXQVR5KesR+8xUUYXcobahdJYf/8q7sliT0l2SGAm8LVj5riyH
Y976oGzCb1pC1nnZa3eCWJ4R36TVU0Oehi43iynx/9VJ/2uJaYB/C42faqjTyVLizM6mK/C7XVbL
hUm6WTuSaVJpnS8ItjfIjkD872mOvynEijXetRfq9VWzKkmYBDzQkVkCvT7nJknK1SLMQiXbQczE
fVbYNco3Rt/DhJvkcjawTolgnjmChsTrH889riLesczqHHI7fjHgrqyebXoYFIhXIls2VIkP6ZpR
aKX5Zrs/EGo74t+6BqVgsvXCbzdeuP+vlb9eiLWakM8rtxPHtIPDjNVNQAokqlqeE6aR3E7LcCZy
8RRCroQ1gX8bbL+e+0dZYso+7I41ox/iDXhSTo3bJAznW+MSXnaOEgOs0IhmqdIjQE+Qch3Bsc/h
LvEu5pM9udh4gpW4grLLYZhjqk+Cz5vlgM+KikihafEDVy5bLx6XN6N8uecPT1JIcCfsbVjQ0WRh
/DzX0MiLSWj5rUk3HgoyDONIrdUxWfLP3qM4Su4BWd55nJ0QasDUN3f5+QcMvu3zzzb+cjqF0YG3
Wd2TRYUHAP0Go5etoBDDHxDY9NEtsXv360CLvUKo74ghofutP4wXpVX7By2E4VF7Rj5OpTNHa3+e
vYf/IBhdbU3UCs7C29tSK3JS04NXmP1MXpczAiknRlXXeJ58dPpF3NntEz6rpEiduSuoNRO+cnOt
22QNGKyb8XRBB2RE1tDPcNWtSiDbR/xTVrNEyTd/8asDZ+9Ke1m0GyL/ic0lMOi4PYy0dPvLHaS2
Kx0kHukMImvIW1RbaE//9UM8cQgit6GiJjFlP00whHZEGGbR3DvzBHjtCsCsUOgjrfrgZrVM4PcI
zr9T6Tzkzz85SFGXs5UD+EdhVyGgBEUPd4Mf5GU/w3IpooEedq0QXqmTdb+gTfUlvjNmIkSnYgcw
4U8Qh0W0TfaqwrYNdARG1B7qGi0wjG46oHwBIb8cMZqJCgvhABI1hmg3fNEdPJelIuGQaJaqKbOW
Am+0KFpFCHoTq4OBoMCvuP1Hp9B9PbYiPPeH89xO5mbS9V6gprrIXWuOU7hMPQuWBW4h7jDPGJuZ
n6RVM9GvXtDi0S11672Bv8X9c6QRM9TsKg3zsWUwCsk+9RfYeo5fpVHTBFahy6gUbnJZ/KEryagg
OJ3FTJ/ps95t3nOVRP+4Vh2cIEJQd0r3PIr75oSwIETj7g6u/YX4IdMYitI19zXiabbAwqqmtFPj
IS5S4zGd1BeCLo0lpbcvW0lFMRyjA0ACy22HcPiHRIytMVtwbr6dKNvUnQkYnJPNBMLVhB5HumRA
sULyKCZzV1mkY+peou1RPq4fwN3I1T4tvSqYlymwVNE2jU2Nc6ek1x6QFeD+PHVbQ1GgVOzsTj8s
PjLN/Z5a8E5PLCGqKmJpD8z3zwyJ3fYOAwGskq15ah+jA5h37DsvrSBqESyg1Tx10C6uAiX1P3zo
WzUs0e2mEQ4Hbu85nY23BT0v/7t6ToZSWWk9YziXi9v7zCD3Jfrct0rb0fTe2s+eqlk4CqFgi0TG
tIVIoqWYLb397XgTyKab9XoDn1GGJOFe86Y56BGVeaBS621Jqq4C2XYV9h9IASKeDL/wDJ4+oEH6
nBPdLwZZtbFgjUiDYdLfZXTfsoDMy56UvBNlFoxhE8TGIYQz0eB1EIaHQes42kMxQtuht5VgV+W4
ZKdUBgHroA1TLq66CiSsyiEbXBbIx85crCXAPGwwml3T4QsehFh0JjYAIFbPSJ6aCkJ4KQsTii5F
4af1Kf57ORRx5ldSSZMUEveJVv2o80UuNphCTtcRrU2nlxL/vm0EyUSKwr1DZNX5LPtGIg7i63U2
xWJdmMo6asQu+TOfnttto09GYOXpWNdHn7hiwS7eiBReKBbiiIG4rgxJNIszz2a6PIBZRG5ozsJv
InXUhojCbBpJxEe6yttsYf0o9YrZJ90jQuI1grw+qiMTlZZuwV9P6o+Q5q3UKnFjKlH+x2ZYaHW1
QcmNWawSQ/xYQi9nDRMiRyuUVa3MrRDctldfzj/dt1McqNkK7NTsoQJbc1eDuPVkgZZjFmEw3CT/
YbFyNz04+Jsl9ZLAEwoRRjQ2XuBMxlr3zwcCFphMfc4k3T1xek/bMEI9CirXajFI72rR0zcOgMOL
kn2qdh4GgrsszokbcQdyVHJsJW4C6cpBHkE6ELPKcxPvvitt1HNuoUBErIDjSQ25SjrgYf27pIpu
uWq6WZMxaxaMW+DZ1vCpCv1NAXHTsnbgA3qbw4F/OY098dWO2OKIvxgpPbPpBVLgS4ifxyMEcrvD
LPMipHYWeDTP92hEhHI4BnrJ0MREkgkgc/qoY5lvn7yi3zzOxVDMWjHslzDoP3/zDr5HM6hznG04
IM1snicWeZUV/oLuwdbxdgxqaB4aB1rnvIMEG6OOiuSfRK6FoyddpGdSJaB0Kd/tQnQSkxoO7dpZ
7c5ztTVhx3PskNzuCrw4GsRACJuI1mbVUkeM+JXqaOBNefjqrB6ZDf3LwQ2Ql49g7PzH2CBnjV68
Fd72U8XKq20YCohqkHuqwc+KzCMutmU9sc8q0btHhS4d51ai593jEw6xD7TNd7VQ9/jJFAcW85ML
ji8O2y0Xqf7WcASHnNj5QPDj+NGVCeqvXtLmZhjkBLls8kDJYv1MlV/odv0llhuegnHHHVQxi63H
in2Xu8cKU6xrFalWPRBxmyVD2VC2zRGSNsA0lP17Qc1aQ/0xAfL8px/icNesVMkIapV9C8fpTtSQ
O5Qwq2D74b98Xv3rMrB+I4tDQDBQpHAvGUqQ+VMh0jkpkU1QDAIrD/mBhLbIpjXIbZ5UKbL36xLS
yMx868LitTkrnOWhI3SDNl2JiutVRRXITqbRDHcGpgV228YDgsQRGQdz92LikHT0SBYOvnXhJAZi
hAqsFOp+xSCeDBO8Zqrwx+M6Yhwi3ABIc6EH8hLnxDfXAovIo0aJuMErwvoqwP9JpUou7i6eWKVy
1UFIuJnf5pr4vTWAncfriacE86bWJMzzsOeyRKvxQZ8U6KY1L72cOHOV0+oyvfAY6o25dwQTe5zD
pi1PkAPT/zBBWUSmRyXghnLEdJZq3teKPjvuZNYHgdDR5/hzM/OxTzNcmU/TS6v4E5FY+fDM8hoR
YcOOxtztg3Su3wtnqTT0T0Ad0Tmj6unK6e+KzFPOxPVppFodmREJOFINmhL1JkBC2GQjjX9MPY2T
REmUV91nu6FLCOhdXV8LQHfata4xZHuGs2jWj5XojhGludyVPJooeLBDp8LeXIYxiwDSbtAZ9Py8
jedIdutOVgavOQvXDAC2LPLsEXANkASyRVNFu4qYGwLyh1IE5xmFUU42e38c7Jilep7fkphHcCkH
4aqqZ+x/xQ9WBx5ugJrI8xCA60N4X19sejjF3VfTJbiDzGAQ29knukQRN9uOPIs9C/A0Esu4pmGc
Nvmsn11ZLwmEV3hz24mSkFVF7shxSTSgFrAWDQ4xcQ0IV/8kUfgpBOvVGFMu6x+lPq5cW7xU/HXz
1xeVbSUHvwR+haAQJJF7Fr2+MXdjJzKAOd4tQvYve2+6mopYkxZE8f7dM/sI734ZDDfUM1gOWBMJ
xE27DpYZtnzQtiVtzHoJJNdGvufKxXnRVLddTv3smdrYw/48hxbbXbQJx34wk8hiX+svHKFjaalG
CieBig8rgV3KKRpIEfsLsgNJx4o6cylFRj6358E5EmPY5goAsAqRXOgtqBp/w8giBoUTIAB3zfWS
FcHmilyDrlhzJqunU9oSqU0iUVgWLGtXoJrKxJJF/HCcb8GckITGyYIOa3H4KkUGPvFKqYkKibkF
otgpu4xn1BvicG80mH2907G1cPnkXZ3sUEobS9m6QXjr1+FIEuHqEvWHtls1y5/Ipfdb3rFKrD8j
QKSHIgly37RPPOGOWiuM5HqGNba3EXLf0oejuhEjlT027uj/tc0GHeeX6LS1MbbGP5tfbeWmuSx/
QPnVWPMZ/UnnAT6C5yReUsCknaNDyZEIIXyziIPR16KifUjhU14YhVQe+U6OtJ8gSBbIyVllv6fq
r1jW5WG7ykMtjZF1+v90jpt6W0agsSjMv/aDZCCE+ukhyclJf+YRUhSeFVvFYFntzqRJ74oks4Js
K16qeaCKH0PCRvG32GE/xSETOhEStNqdWjvmiaOwyWciEamVdtbCfDA6um1XInwSk6T15xEGex9z
ULS3ED01Q2c56vNG1/G6FOZvXPW/GRA4BqVKjtRJ/mzj+JdNax0AHEShYm5ziHe+FEfUC7pMpkRc
Nt6um2CeINrRh4NzOHhWc43jxPbBFlwMPqL2BNxW+3VpOsxpBnNd4jh1q1ZMrAsCC6GlO9hc3Qtu
n4H0Xy82Bq1AzCrw5O6JSSlCA5XFcG0knG9N8kSQSCkm13KF9k6zaHHiSrpX27B+6ySch8fM4dzg
Is+8YjvcVfwt2NnZY9L2+/XGBoiYKKdigO7hkkbfDZfL+4xG2Py+My+bANBbjBxIoJcn78ZxB2s6
XSCzc2cY8IiIwtTIoxuPiO8erBw3S4Q7WG3B1VNdeXdjyNGIvddDMJAMU9+iNy+t4wCiPaffh+hP
tpsdo2RuYSOTGAsWIK1HjFVCDkOECbimSdDklAa5o+nrdmnOEAoyswHHlQbTEo2FacRfiDigqwvO
rblsu+JKVDZe7UDf1fHD5fgkWVrCmquMMhsQiJdlaXWqDvEI1VaieXhE9tZuwYp5QsZRTImOJ/jw
k7IO92fjM9wKPI6YunhC7lefwb5uDsoo1JUOKEdjjT3KrN24mLMFTqbvGxuofSjKjNqP22acGtvQ
o2uPrerCHdP5dZwDRHtCTdfgtYp2thhQN+Hgd1Lzm5YJLIbF42orB/N1RcGJBwd93pcXb5Yg/czT
T889LbQ0t2Tfv9T4oev+kM/EnaVQ2ihZAj38opU3YUO2gxaJv/5xD/KJkpeuAOHGhtcUu0X90iZs
G7tj/7UWgLFUYnDPzZJ4j2oUMa4z7ZENwLXPUDumidBbatjViEnN1+CKRQQccPammFyzIH6hIEdK
ojwNFVWB2ZYQj5JyqkVbMMZAzVqUl0fbYTvaIi0FEDbf8XKBXdeBARE4qLTGfRsoYnDG4HkEvfOv
1JOrYMMnUY7DKZzDelYPW9ehOSaSNWw4MfLQIo/B5HmvJyCdqPUrkQ2UwThQy6m418UwF71iiAd1
oX822YzcaNRlCJMGRyRhG2F6dAV9LCdyfbJqrLhtKDtyDPdjHh4Ir9tlgO8/sza0atOVP9ZvtLjQ
dqjNcAaXEbSHd5rwH8Mjbp/ic6L2egj3ClK+2fzXp1Au/Roj2s/IzE2feeXIyYPCM+khtfL8uinW
/ZM/iloS/8SfaTRPwYWXktYcTP+StuwSE5A180iLXq/hH/be9bGqBBgBhodeusDfhUyahiyXHhSv
CtInwdBIkyMo4TqagGdzQOib/pBNdM9g6YNEN4DDR5pyMA2L6zGPgDNnJYCkzwbirVGeO8QFeLcr
Lv6vTo9CVNiw10p7iCvIwI2fHwvYZcqSwCePKJYrMuicCOE9QBarqzZ7wueOzenT6Kt+Ayq6M9C6
k2EUyMl4A55qW6BGXuFk/XBPxkaPrqjm44K4rMMwa97443BnuKceXQXg5gftWwIdtPx+N4yBpofA
+AaySBr0YD0hNZVo6/pgC3C6dQH/YCnUQiusU0nCZ4PwtrSKRXNwQg/OOGJjnXy3iAos3nGxqaVx
Rl0jNmzNuOLnvAqf21LlyOzJ5lsxTOIjoBEA7xODF8czj3lEK+WYFYZ+Q9FGejkdqb64GRTgBeKy
MfVSIt4Y48z8kpEd0EqV3NXsHQBpCPma4bzwkG+6qTqZt5qYWpLizpbn2VZ9FgqibJy1gutUi9rl
sR2r+HdHO/7zvU4h7euqtjwHOdVogS4nT5YBE0tluf72F8H7lwTE75trFhC5mjwkBuCBRZTYPJvM
8fi1ViIFQtSv8hX6mgoPpqVbwZXBs337zkcL53++LK2cVCywkreMK89ZpUg2lfKl8kuq1clfTlv/
nd280gtkVzUvZNkiKZz5b8iVSsADArbtuMnCo1PiZX8By82j+JpBqE7qjBIIngJywqYfFA6UsEzU
RmShp6XtAhnd/ucwRmZ4FEKZ3uDUQYIjnoJ0KVijpjRV+c8XbL3robH/LrWaHXY9swDvfLo+KwSX
Nd1pWECOVZEmIirkIhzIy3tWHslOzILjzJE4y9PQSYNPFktvW+DwZQLb1CdLIFJZU+dEf1j1Ejrt
g7bsivXQSWkvQz4qEHcMCUJhjLGZ+F8/ypPv7++sHw6qbuk2ewQxnjFbC58dcgDzPvyonRcFQNWk
wI25Q3S94rjDZaNfLdqMBYOlzwzNxrOmstT9Vo1bTS0wUTrZD4O2bXRqAAlgfhqUGaJgPfhueOkU
+fAABk0z6HkncIDrcrUYXesDA2OY5nv0+tPMnWvhLAVZsLaozI4WslBD49oAut2cD0gJQMeAL9C4
N4p444vHh2IjOz+ffqYlKmmVT/fquw5iU9FkLxD3zrcNqb3uvBLAu750S6sVOOeh6ElfChwzfLXT
TaZalJ3464Ao4BdaKA5658mdxNST/U7Xuim/K5HF513tlDwJmu5nDvYoK3MpAFMv4WCFY89kvVQZ
kxYKC0H4XdOQe9Qm+DQoW1OYtKh8M5wip8vUSOatsGjcXCvKMHtFLXo/4ZzMwi4cdam7FlE3fm5A
ZwwK8Vdccx9KHVyrUC4GhX/PdjmC9Vfc0Exd0GzUIKEKJ2DAKwQ8JU7lGRgTuNIUpHzYNjhd9zdv
q9Av6fAutkAWJTEuUyI80jCmVmfmcjlFuuGPX4IaY/l0FBbN68nPThc63zJTYBbJTkfqebC44Uvc
S7KucVfF2OdjlvRt1BC3ZXFxNF4EAaFwo6GN7qbNd8/KZbynHXouVmV4pjmY6KY97TphJUnD1RPP
CCw4FkJ4FydQa86JtPDYoRgjCs0m+q6aiOo7pRPfQNCEVq9kcsy0P092Wr07Sq7XSzcA+iglflwo
GivJMe7wZ78R+aYL1/txNp8GxmCZcX9TcR7SMXlBEiyRqvLBv2iUhZfrhSjW2K8X3yfxtl/jsxMv
GH7rcFARJrXR8A9FxAGLyEc9WuQMrqvQGGtsIbgVOJVuc2QRDgkOwvMpTaW6Bu0cuWGpGLKn8jUn
Br0zk2vfsTIBs2QrPVI03gI4UM3WFovEtrvr7IquKK8O26zZZ087fNduCX1lCCEOO5bWaDUmzvW5
2O2OS4DyL//eDmBeSGUg0g6PsbxBJaVY6dSHM5Bmhc4pnLiKGbRKioznm/9IiE4REPheE0GNVY93
IAFNx9cywwlvBF+QCHyE0DF5+trvUKHw0IHIo08ise3wfAPLj5/puQjyuoWZ+/+PrU2tGI8BCo39
ANMK2UV/Re88roXAXDuTOXidUz0U3I79++u4qBA+ISOStjWI7W2HSCC2ouxfDbRr4RZq6roTvARR
X/DQEUS6IKEyd5aHTyH5p1By0+oaggCIBM6zyMkyQ85nFIlbVVwKzlTZUTAEk1MFUgJghDx3Hquz
d0H0g1ojecCR61oswGOGoaOe4RY/7SAorNsbNU4nXt8JhMqfHDpMaxMUyNMUPizr7RspSmMw42tG
y+w3dc1uFIN0JGt7aRS1uKQHvCYW9pmpFTsQruLuBMlphjnc2QinOdSgNQDTsFJcTJCxxpwYXDGT
jgIlfX+4WKZgsu+Npmaebi39eaQIYKcM+mNSXqG1lS3M7sKnVumsz1vvGDu1Wr8cEMyFwx7eWT2e
6vaaKZETN1Y+oDro/Ac3C60VaHP1dASrQKLvbeVHDPILGClfZyQ9qAG4O9Cs57f57lvxroFTQ75O
KG1XGoifag6M7vnMicNBNkuYcmaiM8ggNPiXZAg6AzuJCJNOIYKqQ5qvWmEPZxXccFWkEDPLpKV1
l1mJgFPNKVke3HvI73dboGglGRbYmb+zsLEE44CwY71+PJDdRf5G2VNDy4riZsJ+8b8OaJw0KztR
x/fe6QeVrd6cAYBST/GO8cboFW+Y3P47EHm+i43pmxht+3nwj9LF8RzNAUIbdW7ye2Sv01XFVaKN
WYSrqAamL4lop4PRjEfz0T/yhuUhOlbNCzVccO+CQwfWjeHTjdrtDrWOldtsu8JPWEUe/lbxPTmF
fKAi+JrP6eFGK+tcqOHCHUqPH7bhSMFay4HsCxOT98hkJVyfw1B/+syzazVzTD/sOFIS9LXC5FKi
NF3vSe3oYRKQmwmj4En9Lq7mYSjpTHEx71sDsRtjpoaIHvpZjZ77aaNP6K/eutq8ETkijRJC0ZOQ
Ynz7tmGINx2ksIuHUWMb+jAJA4i8oGmGqYjoYsT7RNQNbDP0soZS1gzK2aX7X+YZ4IbrGF8p0Tn2
35+3QkWF+DNOuXTVuC7Vd9G8PyiFAGHFceJymBvzmr2Tk4nbKYixHCiOIFPpOJyC7FuZqoehxCOP
H6D6PlGtrY3w4ZVc42FpTWFfUviKXI+sdcADbpP1hD3vCZOf0oWT8hlq50dxruFuo89RobHQad45
q08JPEzI96HU9GPcF4gWwWDKrSg6fyfCoWBjz17RTx5doRpxRgtrcO72x3CWXsgsZYhP+fpbiJ5r
FugkkjTaAmKFQc/YvhEpb+AIqPaG1YqNVuq4cEcubV1YfuA9b0GbSr/oO5iocQR5djmrqzHtgwRi
YH0PEV2KAZ+BwLwLigC/5Yn6/dWEGeIUf22rp9hDDx9zmXJJjYlz4iP3/wO67gxSrT7jE9V3wppn
jo3wB9SBARtLi16KD6b8MBK5tnwNCboL6Lx/AbfLEKkTr5+qZuBMnBydEV0EbWdQJYQwDQABwk2A
4bc+JN31xbBVtsJY5c9vJZijogEUZZAW/3Jf0XXcDI+BVfYfNycQCCvwjcEomgt1Hs8G2lZqTofo
GqjTSvf1lp8nhYxDtbcOAFkC9t2a1v8aN5CCtdUt+ec/nITCvj3BksNW+kYGFPL2r4uNr13MZs3s
vfk4krx3FvsUJxTjpq+80OspZFE/UochrHeu10LUV1q9c4teyu0zBvA1C1YiYK0P5uKus4MGb63G
a4xnJvmQdxyA103WQBZGBq6SB8PwX3mtsoOA0zQRCErUBKi/nyWYsmVRsGnp0g4ga2JdSDwi1esM
44NLeVEujBfVfKLq3NtB8EVXZvheQkK/m+2JcvDZCk9w78UsbjvQ7ljl2q9dWC4fkN527OgzKk/t
3pAg2ZpDssVVYt/EIcKLiya6KbsubuzlYUDIXNt5kBWlZU0SUetGmXyiYuNcXo1AZqybtmXDMlWm
MWnEmu58tznGhMfxQ3xRCMpvtgLXjnhZ/duPCTbjdZ9jiKGFlLDLecfqZ34rKuQiCNLdiL+DVey9
0wAppfepRaV9wLwHbeDCpsAfOgPLqwMcxIT4cZHovdQa0+RaYrcmzaNS/305OGXIh2DZr0NKxliR
HP2yBBMobZ9hdu+05H4MlAeypVmCRf7GDN/mZw+9Nfv4oRWot4BpVeB+0ESjgy7jokUhgpW0lcfD
A7KDt9xJ2lt4ywm5N1S0Ii1HZNUXUn6FFuXPqgK1ADFyVteHlhcfV78jqAZ7gjJ1y3k4xiITduNn
RKZrW52iL1wMwBdiJhbmS1lfWTSwQ4g3bYUZN1mBhb8TkMHm/BZhul1a1OrvZjaapIfLUXXz2UZF
V6SwQOuo6UGZta6yXl3l5Sg0Bc87k1Fiku4/sFW/MvjYIYdFJO+KCpGigsDfegYlWCMH7Z4cvi/D
ApQ+9fa6MN5vjjndrb7YTupNYY7bfrt29r93EpcN0+VBYvFlomePx3Pm6U26PcKBC4f7P3mfFrYE
NPtPTw2eq952LDs06OjEkFofMZYJXZry0lodeItx1z8/BtEcTrBykN3M+Ex8dBxxBNpV2r7YzV4l
aR4HivSF0+1wA2CnuAmxIhMcA4531ecnhmAN3bkPVYc/r9855YSCApA6C9Xh90TI/6cAWx/IZSu2
u9humoUZyw/s/ZeapDlz/An9lo8Dc6nW0Pe8xpgPZ7AjmWORgfGBwXpyPQY/VIijZiLeeJTQd9Jy
g1tqA5tdoPjt9hUqN8ScZawemn6EEDXQ7erIC7DK2RPStxHm8h6Ivb6/KYDNdr4wJSskGrEZIWKV
PNkFxgGP+zNdUdlVUaWk4oH6wB3+lODSzCUhwrQKBzgH2brrxHRBkDNH2f2D6ImbsrtAi/bU3QO6
rUYQekMGo5bP0mnZetQyU7nustgtYCxayocD+z6KWKTLbr14iU+4NGMz91asWUZh4oUdw8v258w2
a5Fw0z3b0ItAOnOYnxp/PjdWHnGkj+ABJFFbDSjz/ZoEMoTvlxpXpXG6FRVea5P9xMs5aWyAnI+N
Gfv3WI5udoWke6mLnACUU+JYy49KQlmYfC2BZkLgksfK1JZAsvwpOH5lY5yn7DrBZOEJsUWL7uk7
0yZUxt/YoiBNl/E25IBM7RBuQE4HAOEJDSh+F5kY+CPAWuWLgjceV2Z572PVv5O+meFIQf1pURP5
1OjQ9DqTkGcy1SPzqMg2Z4kkZrnLE0S956qc4ymBtvBva76+G4vBLfen1d5CjoELHSe7dAue3IBH
DIAEI5WCpzVGdRcf1HJeGO1crsrwH0PLVRuzjfTz1JMJxBAyrXQnl+49WjSqaOGe9Oxq3MqqPyER
c7y9Dmj1k+rfZXoV0LhOQ9Baebozs0sdq9Z7is2/OuuX7WlqdK+AqIlYsfVDbp1h89PgXMOYu543
A37Jbw0FMvndZwpYfYAb9P8LRLVWk/NeZcrA7+qDai02QwNitLOEpxMh1PmMNpmdLcR3ZwrdSXyl
bhj6VckN4wRXvelsZKTktdQ/C/AzdGQFzHKXj8LriULfsr15rOSvgFThaQpr51yNUX4qu8X0+Sfr
cB7uShaghKE/bZ3BQ233FctU/OvhHiJxG58qnMjGbR5gL5SA3j/R2XLASftQ3xxPFTmxtRBJM0yP
KfkpQR1vzmS+Z28oIAFtjOnNCeYtdk7FUf2NjYLHYpBlJF/m0OHAgwxbQGzkej4RdlE+TO6wkyQs
kCp+DjSEuP+VpNDdMljjgrtuOHCqB7vqEzZ8GGtPCVTtyk8T7qQadSw8i6F6bRi08rgroo6pCa6v
ZsqwKTu8WaUza64seUoLpw2vwhGBwz7NIIE6YC+NWY6Qjne6Jvx6LMR3PZNj6VSBOog4DBLC793B
sgvs92SqgkeZhXW5OzEq6MR4Phc6GY0dfxUD58UwrY0hLlh9i/hmqS1/tfRP6em+NyR2s3jbfeOd
QJFGYrOUlj9aXuPIs8BkZLar2yCe2gK66/Ylw3P5UB3KupJ5Ick12u82vzdo6c0mNW5bJIH+NrA6
bUG4/kPL/oT8jjHt4SviYtfuc3UOuonQhpndPll4Z3l2e6Obyc40hzbNqiPfBN5mrX5eGwNe92T4
OnX3cZi4dQ1uP6PDdddpowHxuP70ZsDT7m2kPuE/IGO+M049DSoNK1P/1v57XoFs1wlF+bVRRJeK
v5NydeDRFpN951TdKsm5y57EieHbtSOiOhgbUI21vvIDoHm3xnCInalNED2koe7ms+mBTYvybbX5
c/dIapcC7yTOhqI/HMACzHSyp73mpBbD0YK+mbGYur12GB8ixiW/YYS3G4b2TUmPnulCiQEqNhHh
yFLUL0UDP4ThmG2EY3xcdoe0YbE7QBFXOZIJkGwkiK6gzDB3nOsB7oLrYywXjnaRlzPz7uPtbd9n
ITfXBR2UZuAaTfhGPds5uYe1HnIge8dD4GvUx9hv7d4kgvSD92W1Vey2wjqyUXD7nkYEvuJlNuWF
98j50FVYIFHQzGIs57RsnTNZZogF1LOfUVG6Wjzq9JnSeyumHu1qFKKFLqf+bCdim7cYSKEvjTlE
l6YFvhlnLuHZ3V0ohq+pmbTOF/TzneRW9GATDAPkKgQLxThkyzaEEau8M/QEElmLXuceq5Fb3vmG
poZy6Ejj1LvzQF/QwvkveY9OmR7zDXtQ4ZYKHwhE6Ni05vzkmA7GV1c8EgeuJi+AHdVitHrAmdrH
sadfp5m90pxiaqFORHHuR4jtkZy1mDCON8fA69pPgv2zXrlPSvM9SGf//HH5M38NtRS/1SQ3SmoS
BHBmaVjShz6LZGkCAsD8MaZR5Hy6XiqvyuTaNRxsb6o+Kuxst1lyTEm4iDabqvbj2dXCrc7zg07N
KvWgFQgSxZeRjrNU6CqVjl9b2rh/N8FlXP9U6ClX5pLq24rpuGY6R02ruL/nxG9QRX5QhOzyoun/
Ajt2DBAGl9KbMBQSat9/WwTM17xMVSbSSSjqVdULR8jqJ7teF/kcUb3jwpvIkgYfzeMWlhu3rc8u
T834/SZ+CXoEoJQvGiwsgTwDtaiqpF0pQPwpNh3a4KiHVnnMQNS/80qTfQfVdxCUkr4UA5sHO183
H/rbRvGzdgdlcoWFtdGwvHRoqMEQqHpdGPByNypj6Jrz87DgJNeWNuIREIIFlwmyXbHrEJJjOHvk
7dZYMXBKoF/gi3W4trJ0yT72H4ntaS6wsLil/uR4X1FADuWpj/hw1yDn9hGXcnamY944kSlofTxS
D4lIeDkpknViXdxqAFhAQ6DsC5TlCCgriJ2VDA5ttudYfP7hyTpkMKm69WGauMSqc76PgPkg1cm5
jG3FqEVNqt3aNBj60tuN74ZdwndHpy6lmEpQer8fels/B503JAjoS7l5r6yAMg1RmbYdz7ymfl9f
sTHFdv1m3kHzdEITypCXqJrkTDHnFTBBodGtpcHl1HQ+9hldHh3xIpTioDTqendtwjyfSWaAs2Dj
R0PxI2USNSV1P7nIyiJOFzkCWu2GMmMOiS0c8mAgi+Dh0kljiXdNIfIvCez8VcwfgDigqEb7YKwB
yEY+q50XEfmswPBI7zN92L19VqPzokILOkLZxooGcmeWj8yjJRT9Vv0NaKrMoxs365SsFK9Jr1T7
kBjbO45IOtrdmQGSVVA9ZgP23wRHbECdgPoUFUDd/8SnzMd3hONcdAa1TFBp1flACiVjDhQuOIV8
8Fxk/MbQ8syxI1gR2RS2k8F3e7SA06E5ikz7fxUPJUk71TX/0OYvj5xBIBX1s7yUU/dnCo5F8lph
YLExdWSkWp6UU4Sfcb8ztuh6c2qo9vAzHSXIFAA6irtxzgyiS6YGCZ119uJm1okIWkEmz19TGQOe
UNQIQUwDBsO6o8UiN2D7frqsLO/MePJToKDzp+tjj8FLjh7KxBUUOCrufQO4UFCBVe/AVYqqg0eb
MkrYEOkZVjGizv4pahumdvQh5g7uQApcq7kQfyItiTc8k2cXWutyPaBRwRSzdnNsHTP/ltpDNnEj
RB1FI8cNsqjP//8OcIz+i8698l0T6pLZV2cucKE97OrXzUASG9gF5gVFZnvAVmvqXO6kpa4iLyJS
P7ZA5zt84wwpDu/Tv+pBZf0o9zNuuGfB8csGdO6Uc0toZp+wt/aBVE3yzr9tqpTdI/I9OasODUhb
elQwpSPy12hXg2gqKk10T9LwBXZ7kIJ7joJc7FEDzQm6TvzoiVwc0WC7EOIlYT+bkN2P1MPlFMjw
SIEazTH827SoUYT9TudAPVbxlsIZsgGfbYk1nGUIKAe4SJtYTKnGexItTHlYs35ptNrjFCrZ4OYM
//9jEQWwdJ5umGJrPKUnXTXp0S4UFvxAaV4J3RzrwkbWLz6mS3uPlO20Op3O/nAOHp2SMDaugVka
SiE2zEkblESVTEc+DL1gx2Xyia+MRGgYV5wEKsoqkXNLexhpzNb0+y4Bzj+q7bOdv+uDXJ6vbZAY
G4jl5bHXKjs8vGk/Ps+zcy490ZHZcxSf3SygKi6zmd8moJlTCKtz5bU+4uJztLsjB1f7cmfCHFOR
ObFzOVNRnXrxJJREVCSClJXFEV5RwSztRdCJXVg99FmACYacE7y2ZMojmICQuo631c1tn4r7GbTz
2zPdUGmUf77fbi1PG+ignlRqtZgISrPR+267hJ4Vvefm7PZcMboBi30OzM02673cLjByvdHwDceA
uvwOzcWJ86yLlt2i0rFIBZO7q8V2JxS+1IK/CyZusQr12CUIuyVcmAZ8npfkmE7lyRQ+aV30T7WB
987+wpGnx4cmxpu6acojzCsVVeU1pJSZDE8kgW0427DwEh/1hBmQkfWDfd1xrwXDMK4BBSn+6Fkg
sTDdA+HehevRXslczgEeI9ZNA/dShiZXhzYyoxbXvacH9H9Omz1+wBFSRcsBJQJAunxbIFDmlAmK
FjZuZX4Yc2OnBGP8MhT7LxgGTuIXEncxfmfPRQpI25nPEL07Ji2NhyyGpPU3DtvkxpS1wlpwB3+W
pXB0sVxr08JvZjktLfMUSIe9oRfSnJbMZuzFhANC9ou+bTGwBwmLF+RT/PKggZygO6vJ+a0UqXsD
joNSFQAqIUbjy8Coh+JWs37kEIYqJT3gcr60HQ4i7TqqFVu0l0sL8UkXg6T4N2IqrnzML+kptIKa
WhzAxtO4d84SyghVilCN8QTRGlVoi9G2Fv3Wu/1bjf1hYAbLB5pJiaeesQ08Ojdk1wtVJnCy1dfa
lrL7mb9LPbOo3jBW/pWtjuWSPVkvasARYb98RHtO74aIXgcTZGufxzBKnPh3q05CdS9YfNeQEBTF
pIr2f3fdxR/rKnFWtDm1GeV8616JulXhet1yliEqyo44ALS8XPNAvfZI4NTZb5ATtga+MxW0xdmA
AgcJ1US8MsUDuUY+Ro7uKrsw9q+jLa9/Nxn0FchnFGd8fNI8hDAUpSU5ffsIdiKYAHLq1zKJDalk
AIgsL2fgKqmmR+bwbKh3T1jbLxL35ahYibN4LOqTHK6nB19k0qvZs5qb6hgjkvXNea3HY2af8Li0
9ii6eDqefx0apzJUWr5OWDh1LkEPScA958e/f4MSJNawdKq8wjZrv0JeaE1idKEMDcKXyC+qRrAJ
8FSl10+LRnAxMK4Ln0lyRDs9tU84YNlG598mSbiq2dfMGeaiWAp9TM05gJ3OpNokGJ1fbtCMxysD
YEsvx7F0KkQOFMsJ77UtwU8dei3HA96hK6I+O8LDXenvg55emCaWjy8L8USubt1ozsWonrDfOMx4
KT3dCCbMTW4sOJg68cvJwicevIxeq+IOxUB7IJnKvifm3NFRwGDoAZtByFfu2o/hD+N4PPnB/uLb
ImVDyQ5JsuzyBuCzAKZ2KoaWhAgVbuIq8zCKL6E0Wr6pXl8ONNpNkcZnxlE2RRJHQT8IO+eWRQMj
nldVUbbZ2sF+2AP07lWah5Q40S+gKSI50PiSgZ/+q5zyCg/RSSjvTtJnXTn9Ik+F6B0juAOb4rEY
KXSup850qY00p7kN+zpx/zUyqNDGE4hx1aNHVoCBD01zLY2unqoodKhszh0DlW46kWIaGN16uQDV
gXtW4NMs7SpMlHAQN1ceaAUJhPAu7zAvbRDUFUFj88XpCIwTApabpltjLpiXHNJoDn/i4RN5YhHd
mYR98dei3KtqvCGTy9MyJn3iREfBjXNAKnK59eEgtQoJG8HScSPIQ0Gu/wDHWlkMYN4R0vLLY92i
A6NOKLHXETu17VJUmubDFZucI89cMchsIKzWUJWUlpnY/vX7OnC89PcoUA5KIj+Qd/pQ/s6pL+Wf
hNJ3E8w3pqF2nnB+eZaLpgB6kymWI0a2KBzMzKyTLwjxOMo4YHj9g7KhHuFh9NxNJer09sSLQK1x
n8chklKJfxzzv1pGMc89cKr6qG/aAg3cMHWMUz87RfrZ2DXIaC1tevyvMpNjb/a6pqJaYNEcBSGo
pCB8Z0tvZK9MP9BIfl+oHi8TLmu2JnKhsLwCVr0QShnfduZOIk+h2AX0XRsEkk6bHRENFP61UCx+
E7hg6c8g4xSE6GChNLVWs1WLMGBVGfw2SQ1tAQjkVC+oIeH2lmh7VS44GNuS8EhJ2szarFJm3Iy8
sQ4liPNPqR3JnhX2Uslpn3lNYIkaX2yf/zHDNjK4ChjUIsp2tAE4tL/vVUW52Fc9HSZcfOhXGXWl
cl3fh48aDIKzr48Q4FH/YHpochNgGKdzICKKtD4P8Z+FneGqFte8TL+Rk/9f7ua57Hv25+IRWSbM
LIzCjIgQ7eMZ2y+9zCW5wZUojmxF/TaWIyoyDEMsgAPo24Csd0i+ct3KAd071Hm/NJ3qfJJk+Q8q
zmwFrQU6ydIvyh0MibEUfUtAYjmDXjNMy/jp4I+TPfHYvZhiWvLPCuVWrAGmfHCf+c5L3uHz9Hmw
peRX/3vUFSSobhPSg/BhaejQY/zuifcr/tbajaHzEO3Gb2OvWHqdIW76EejvDfRbm5TnDfpxb7W9
nwXhWHPJZM6Il9ijJdgeiUHUNEpvH9y1MxdFhnhNdQ7haVKFv9ao3OoX3NGTQl4zLDim8jd4i2GG
Y+kbqHWo8rkKuXxaXCRMuVxts1FnEpa1BgwxZs5KDoYxPu3dt0P3T6IhOm3m/h98/m278pe4UKMm
m69HXwnLvOEDPrE+7oELIfIjLf+ow/7kFau1Qj7QAF1eWtohTapHXEUmn34p491K1XhC/TdvVLpC
lioc8SUYYj78wRkRezYUykfYtAKokjykkHcOV3SBnnL6idsApOePsH9T1YoPTdYfOhyKsZAnlzRE
t/A8Spby0tULOvb6+Fu8BGBAt9j0dpFMHDpeil350aXb7FbgwLmfqNRPzAKMU0XI625HzAIVLxLT
34gGuSDR6PYvS7OpnygTs9AznR5oDKZZGoRtfRN/woMievePgkxr323SN18S+yhyiLGs4QCcBJKC
KttiPhrAGLGZjbTZUmCa8iSK188icnXpBZolq+KX8FmDMictcEyXB5kZ9U1I8eEk7uPZsPXd09Wr
KEfT5xZU/HaNeeWBW4S33dyP17qRTFi4EINmfj4enQFztEJ2cVgtTNE/mPYts8Y2k+At6nxIFAw6
Rhu9Yqh07xcCCxDZ5MfZONSh34OCKL0ggUobGHwuHB9h1SM3XeTUmPRpvCPxG72t3H+o2DNKCrlP
KWYzQawMZdYwX2PmkWaaC3Dpf99SB9LR3p8VXJDUH99x6ouuiFEHOIQyXyvRsFg9OuJDlF3YJyew
GCVDuOmsoCnjVy+Yd3dELkdXL+KuVJmqTS3k+WTkjVLViVkYpC6TbidDj2r26qqduhpS4z5dAxIL
nAU8AEFofV468g9XTJtmRP0QO1AE1T2XHp7hmVE50JlpvKiozsNve4JzzIH3ZCLf5z/I3hDydRaf
Md9cNdQ4320EKlGo8tLz+LaeiXHtt/nD9n8abwyWKDsssqqB17GNi1rZNaJv4VgW7WZA7XB8o2bA
hH+MYPJOUMzz6qfx/WDg1IfL7oBjO5YJ1pyelQzL66XoRfosRprQRUgu4cY4f8CQCHGMXfSeNzBO
TR7JsenBZh7b/aUYcXZ4PtI7eqssq50fhI8dvuCwFhqrNnOGHAy7pNcmJhGwfY3z5JqZV4USLH8P
B5XhEyidrYkW6kT9H6xiGxBbC1KDZNIvJsq3EgpWbxW3M7qNEynzJC4t9nh/NEIy2OJ1XQ0AirjZ
oxqyCPCdPFH9zY7DTyUPwaoT6W65iWsnM3mFggf0VUACyGRuXwjpuvf3tLZxe1OtfKvw7ckjOOrr
FH0MBs4DK71R6zj2CXfpbsNoaJe2HtKJpj6GtLGbh9CaO4dMF7QIAdUyIDCA1aHSvsupBP6ZPOxL
flR34Eh5eKCaE0V9eL+i3o2gb5qEvzI3tzZfvIpePw/av7AHv5RbQ4/0dtDnFvhoXYdNGxppPKGc
Bi6bcWcoaY+0uFdqIAq2+nN5mVgFtW1JUVB0K+jvqlL15ythhcHghSVTj+TpEEY2NgILZohQ6W4y
3BD6SG1C9Ry+DrbaF6o5H/4hlaoK3uzpR1PvCioygM8iIAU/JNNNP2YBHpxNqtWXi0AujkLuWpxE
hFa/tyZUMnWlo/9NfXq/D0oXjKOGUFHG8Pgjy4qXS6qBMOD6iDqv5QA0wL2g/TpKQQfjLcohAriv
NMnmfOIkpdbtjtlNLKwQWsfcRAnVuOOXBduK7TBO+1h9zdh5ngGN3zEWnU8w/kigC1RqeJgsJcBW
gnIAk0jpWvis1ki4bmC++/xgFQ/cG9gug3xwuNpcL6vNDen6kxKNoC/O1Yvar+dP05Q2Rek+KnLT
jtmAoK8fzVv2jaG54h2r8auh9LIR+t9syZxc0sS46sDxAg3YFzkfpX5CKa1wqL6HS1owYaFuCI+C
6EAh2NkAlWO4dm8m8f3+6P5VWZCupCafjTWOaTxPvykWNd1vELTVBCAa41YdvBfK+VZkJYg76owG
8ZDJJqtgI9EzRKidPUzPrTQUJn13MWJmBRNrWTI7R0Tc/qrIzYGuExAvgwO/42VH6Aaj8fW5ib5k
ijpdXUpdT9eDotKG2e5abh7esjbgKcQ712k95m1ctdJVJ4e8I0oSbyal0GF0h/QC1gCNVUI+bJJt
kYnizzY8uAljuFi+MRwNX0oxQ9VTkOQR2o3B9cdS0/RESQBDkG7h1dck5j9WWNT0rcTvv2GmJQpL
f5zcN2rERz65qAsf2MZU7sM9+1wU/QOMFWA3pu+xG+xMaFQwOcZq6AzlPHBaHNSzNB22++xR3e2P
rPaiaKki47VqSYpFTLqpP6/g7ZkC4/rJP9/vINpdASb9v+3Q8Y8mmtMrC/h2IUFIZZ263Vdl8CYH
nDZfgfF5AY/i9uFupevVmCxjohCGDJsFCImLHClQgAyKF3pcCUEUemiQF+KDwEJItp7bjDtP6RGw
GssAfN7vzMXBLIWi4LFGRA69GoCcE1WZ5/U/CYkJtNCmLJ/2yBYRvhk8riL++zE6+0iWce/mICPL
t0J5GyIE601XaNkL4Ma0hfx6lw0qD5rcTvEYzARDz5cVa71uCgnUL1z1+0lyn6UwjEe47FlTzm0K
XogADh2teedfaLnhh0lOYJb0JHR1t7l5yOP20LXZq6gxXgPvZdBQ5P1B+HzUF6uqMDU/2FEv/hGx
WAwcwAzf6zbBh0HZb0pn/6qvocACmT+66bj9Ep2w7T/FwKqi4S3Jw+E8efSVGbPOeu1coad9OzmR
y3AojUg8Q+DC3p2W0vuzmpi5JKOMI/uAsB3A3qbONAyFeraXBN+IZDdn0OcrkiW9f/H6qqUMX64A
SnXg0/Qm67unv62V2IQbhvnM8IzjCpf7kAnSsqZ/j9HGi2N+9ukVCyjbo1lw+hOds4cEUhuYYiq6
gX9wmAjI4uZWtG81yNn8gMjwGnjfdmvxmyLnfugy2I5DUk3fdS9ojKkaGnxrJXrugZsCzWIc0eVD
jmy2iQSg5TeyBIsLBkKN8tGF0dgFCuabZhzKKSxcOhXvSv/bPGmvRu7+HMfOVtWVzi/Z99n1VPhn
alpjeHfAc1oHs1uyofl/JPMk8SAlRjipWqnDWtgP55erC5xY7L7Om/MJ5njtwzhRfHfBUbvau1ff
HXyh6WvPzPESJkq5Bg6OUiL5ENFsZXm8B1QIOL0vP5ABTnuQgLNdLW3K6XeYioTk+lgKz1U3WBPo
tcaivxY+kIuuF6D5PlblL5UsGAL8/Wh23ygj4LZO2EVWrAlpzzRmWvKdj6AEXNx/ilQqVGSghoPx
mRShAmwG3+VaesD1wvJpD/tInfJKRuXUNiLrcnzzqAHXCwH66axjggZs9NnPIfD1wtKOGSHMBRIA
y3QUqP9+MA1mdAKTd7zOrjHnDErAT+0PAcF7+CucjweQTNwyEF1/QqU5rGK/llApkMkdbgxVofdj
B7qC0oYxvPPGPmGbJslrrp82bpXxN//aoDXS43DkehwOom9/bj82nHzZfQBJXi1R7cEYOd7J7u6r
btqlgQDycgkTWA54Plu6n+iJzDuHCfvuV3zTy6gf1GrMg8p0UaqEyK43iMIbgyF9ID0/Kb4fCBd1
Om0n8KDhmccfeBsWxyJjxJwJdR+nAIBg4K43xk1e+B+ON61mcNrmPdyju0SBxN5cQdVrWrdx/QLn
tmFNkPB3FfMvqTSQSvn/A6G4wtkmOmHDNJTXmYSI1LlEaJaddgquxNnt2H0Vlpi3VLZDxFz68ce5
TMD+HgBFjBCArFIWi3wIXSuV5XY1Lt/G59Rj6oLkg5hY+/EJOlrx5ZaS+e/nvfKdKlvgJxejeJua
p4WnBY23pzSDZ0RhxJd7PnueqfNV+GLigxqjEpcBrxE4a8Luw0GseUntn+1eEAaDreIMN4kw+iDx
nIOEJPKZ8HUb6wgkg1XMb4NFLHyGFIicQ/P9G7uF3UnWI3wFn3RyuqOwJ49A+cT8kB3JAANShjSm
1RPquloxt04SR/d42kQEAqhVhxXcbfY0s2qIiVYmqWxVYKna5qnMA2z8NrcQgtx9dEy9WVOzby/7
37bjfJXr9jboVViDqy4qJ9aTYicCFO5VPvEacZEpKwR5Tz1dBXmTOUjYpIaPmc1O+DF9yKGJaTgL
QqgVJoPX2ZOmaJwhs7zqX9DIGKgcCio6nxYYxVvkBJ+Lp+GaWNrhtwtZZf7kmOgnyllQnNhbJSe1
SEveyeuyY1wT1dSW+QF/XoHNc3si5Mkz5w8AdfXfoGvnmU9xDxG2Zo3PmTReXL3J6y5GD8bN23Y5
Eh67dydesO+mUV53QhD/TQ3xpqilJwpV1x4Epvlm/nQX6axvFaWW+v4a8Q7CxxL4JE+N0k2bOuGN
RJGAn8GLYGRaO5hrM8SJO5zk9aSwuzAZwBsNdNE6cCF18tAN8ykXyvpMePmV7lbMUfdZb4+PhXBx
3DA7d1ijVmkN3Zp1XvR5w9/x61y03vihrDBGt7DvhgkYpUc0dsja/L5moyY+vVC2qtkFw8m/YRhV
+yqu3T6rq3jF0puFzNzG6fMmuedlM40ib3wsHgHkYsVFIKL7rq8aps3b0r86n1mzEtneXuWyeWDp
9jc5GIYRHo789xzWxALAF+ia+CEI8qHTZV+fRpryq/fg9hex1DXzgaE0E1trw28rRDjmnN7rUk9D
y1FPW4uWAu7IsT5f/yMvhTTsG0C+flm9ZPpmwXTBqF4sKpuL5n7mV7F9HIsZdWJHjNXtY2BpMvwy
d4Q6qqtb5ij6EEMlBSa7ZIQ4ajoTWQQBT/ohKeEkiQeLvLKAjKzDiPejXRW1oGGhIPJ0xaGXCu8x
Y+g2hcczLq76DJ1KhujfbsoOy0wmEgYJckhe8LDhl5ulOi2NJnv5+4PEy9EXXevDGp4dHWXw73/X
SEPIodflAUL4WifQMM0k5lsoBxeN6FNGTmoDhDrvGw7erNT9uJUUMpoj8t9hCtZaCGrTulqTCMsE
BQ97aMeuzhNMeXYcNpaUgyV+ldgkFrBBHZ0zXGcw5gLo5Cjpx41xfqN45yIGqHxewcRpxbS0l1QV
QAZ662vlUsSUFjHrYzV71soEs+4AWxNQAndkR2N97JtpTw/yJe4cAdj67boe1VcfZsK6nYeAgJFz
fA03ADo1SoUzKpk7tq5atIEAycvukh9gXdRpGt7OwlbuwuyyI/q6vj3XW1m53CDMTc5auI5aCjQF
+BmZ4PDuRtSjZ1GXIJlCufBJ8u4lqnxzJCa483elQ8ycSlcTcmExngwYkp41pucV72muKkK1hPpM
BLZIoMv0JeePcS9mPSad+9631WOTKozFUfgqUYb5u9OHx0bsqM13KS6uNpa1gxOxszvRcig5OBQo
hQiwrORGNehmv1awbkmNZtPBLHFHyPNzWE8o+zjRkF70/lMN5N+lw9j9v273YgdOL0Hx3hAgcJ5D
74wjuPPA0HsRU+d2wdw7m1fIS+qUqpXPKnuNmHPcUSQzd/oRQDQcdJRLrDFOgJ4epWjs+LKii4wA
Yo1zwN8B3iQavu8HNXOTglk50K81Mu/ndeHxP+b4Ryue6UuTR4IjkLOlc9oJTE6Iv2WHt249miqA
ms0Ej92KgsLge4btD4ZtRb9H6ym98Cu0py1aH0cysWq3jT4H0BDTjsYskcHhFHNC9WM/lLa6X9Fw
qdyJ1RH5QWVKQK6MvufQkFl9pZ+RHr7wv0G413MWUJ8ay1R4OuIEv/w+loQDaoMnXQKXfA8J9P+q
lqfPwZQ0r3RFsPGTHX1fxuKi1qt5rt6WtN6TZ6cvz8fXIShvBZhSHKIOy2SvmmhoVGi0mpS1aai/
qMEBOsEZJzUb6qbclxx/T4pLff3N5lXqjOwQqFeIZKVmKabpKTFr4y2aCVJ93zgz24MYdDQi80DL
wb4OqCXGiBeVUPdcLlwrbKnMU8rIHlED6ygzkG6/OzLS/FQLCCm5w4HfviYbzUWuZCzwx50hJsk6
1ZbcmvYKMAqMKVNxyLYa39oSKcaT04ZJy+qXXBd2uW6rXwKKvsYoPp7i8aujAY4iEep1C2VV2NGn
BKGhOQ86qgNd8rQ9OcgWV7Aw3BOh80buEjLEQZG5Dhhd6auC/JBhRepEuiAIfkCMkzDjynNzW6bp
XX5/X8X+JmUMt9R7XIOftAa25NrBrDhL5A+swDbLvoqLqXxmGezgODAgMhFXE7/C9Yrzd9j64XZY
jX/lxW6gPzRLGjssnTNW8+veF8XAEan6TZeSDgcdpIZ3q/0r2AITzuzSxABliMwysO/YACIZ8Mar
z27qIHc0w9Mi3pEuPw1+CnPsLOJSNc+fCuaByOPiWQ9Te+KeUHb7l4F8vhp0zP/4RdBuMsnkTMXf
HOWkNX6+VXvjHs1mmMi1gYPX4YIIl4dnbxAX6YRKsduLJtmqFg6Xz8cyGG4uQnOGVvr9H9FZAOwZ
J8nEY2dW9aSx/fkRpN9R08r0zD6jJ3sf2p8+z6dPryLIvKfPrnvunZVujDD9CySK7oION8+8kKjw
io0MBJnKrmo2E7h4GzMM/7YOBzO5+cl8Th43rpBVk5kSMUyWUgytqYoZm7GLaDcSjmkL1e9+5h6d
OFCxmWwYs1iOma9jwBJQZepc7kDODpPjw//8cbVgvdopKUIVYN7rRPKJ9JX40gvqOXTFiAuV+XUh
fNuOl0U+3NbLX1HXPDGOp6pePURT2W2TCNBp2529WHKvulpAxWRumreNlS1IHVNdyEMZsp4rlXCq
svnadIz19KeLouQWoNCbJgZTE7+a4Pc7XahxlUD4dGH7mkYaHfddsl+EpwmDyJ7yoisYsdzst6V8
Zz2MycfNVq8BSigJlCegtZT094dz3cn+fPaHDD65285mWgWyitFlp7pdMN4+t65sndKM2lsqskrH
OvrzmTP/QcR/Plk7KGhVrKby+HptfxtiWSSpR6f2ov6jCW0Ml+8Aw37Awis9RmmHTD5phF7ruqb1
hjOk0Ejjqms5RjFIKuU1yCKkTMIzWBSZKYWaP3sNP5aYyKayqaQHsji9YcW9KE6/mpp6fZ9lXvTw
AgrcM33tTxwR+q5EjWtkVpfkjdYvEegshTq6vIzlJMD8slG7KSRsLZYOqQ/YB2ZgYhDcuykB+W5x
Cev4kzd/ztxBAesgWyICQ8c1s2Oz6nNY3Ef1tO5gQKiT5D/9gKsyQI9ejyyujWoo5LgPBC8c+QFD
z4LJxm3GALmyh1qfJ/eTFlCHpGnlhdk7eyfYhMQOdSK1uppQQpLhpHu/+SjFhbL/VzAZvTWWvcfc
wGT7aCPpLeICImmBkDR1gPHZN4ri/aaHKT1hgqJpkLIcK+02epflaK2r4rGsNgd/uI51+ZJnMU7n
K6K/1Nr8oyfHToz8P8Cc2FSFsaqMKiU7RbzTd+PkuOftJgcGx21uLoRqwds1SJkwkI1iie49FpLk
sZ2pX1nSQ1FZF1bDGFV8SgHyyuZhQrPDF7wGOLXlZwfb3q4SQ7+MFxy51TyOrKMN3vZS9moygTvv
L85FDeXPBnLNHs1y4idObaIgYP1swMi/Ua67HT9Ve7x6CFMeuYTJxieMZ7409elrXr+GnGvvecO6
hifIY/+78aH1AXyrd7/EGsbqY8TqmI1OFiHwnDXyfjrGz9753e8E8+FsSkjtJet9iaLx+hUDB2XD
cKm0eIVzgS7ME1FaV8KetIuZzFQbPZ1HABanK4sz9WyxkyzVIJQ+P/ziJdT70rAmE3HQBxxpQmaP
JuBZ8IvvKmXoPOhfHSrPyDxJwC9+9dnYeMJITGAFZ09i3D7ACwIboTE1RjMZ0YX3jylTycXkOslw
MdIr0mcJPSzVRMcHz10ex4z0FQC3OQ6Yp6ZHPP8jfzKm+DBTGNReDCY+Jz4AyBtDSMIpaNxKDSMo
P87JgUQj78zHKPxJBAbc/AYk4rac/maghpeY51s2Ue6+auNqwNsaIBLx24GDAsYWDbW/3vdJ0Yp0
z0GycFWeMAk/lmvyDEh0cTkUjef3M+EHDeGXMzTlWUsW3TIPOf/ArYUwFExACiHQp5Fo4tTEFl/F
s4/814IWpChmzRQH5UM/4Wcj3Uq+vnGBv0PwDcirv5Wkq049rNpr4cn3Yfq69F9bJRaq855ndciq
iIALXKzhav2+UAV0QSXO8/JE+HoqCVoqU+qaosr05kJmQhm/nIUZkBaQbMMCsuHhNvFI02hSANg7
M+6TV5uoYV9APKzzSXfC+N0orl1y56gXIz61Hi9qNtxWh9g6usnGrSKs+5pimDKqznaU9PZpGFwd
7qVeqJrJGfm1Mt+WL5GUKgYu434GVDmB/nDn+2JyZrT0iQ6KJoG6HFP3pN3wljXieYbfzuJY1Rz4
132zfJs3GoN9zeD20k53zY3gP82t/rR+GHODjV4a4dG7Nyh2QBVV2NAGQO4o7kYyYXH0wOwCRhE2
zBEt7RC1c+MjgplEToXgK/NgyJPAmNdmflt5TD4kRhPKQ15MvDyiF+Yx0eIScP4H+TpI5d09V6IM
/SrmxULCnXex+3GC0MiqveE8a0AW3Knj3ry/pJljvccuA/RWC7cL0m9+/DVrX3omQYDS+sgCbrXN
uOYTGwL4fcCMKFhrCIDTQEpAMaASSvWpn3m+QiW1KeQyNHr1kL4oaCefTOMx6aW6B1ufqTLqLYjw
LxxQbwzuokazFbmQqRuCvua6e3NM3DNA7hvhKYc0I46wFZFfFQbciLbzOV097StJlAVMm9DvwYtp
1uZRUwZUxAwrwV9GxgKdY0W0+ltWqsD2m5rKaBRAZj+8yxNlngpj5GcConaZzbc/eUdCvf9R/5YF
OwV0v/0lt1O6/5d6oob4cPsuwjbLJDZ0Jq9tMYsWYjzilRYtlK/vtP9b0ZJIaZPQBr7h6lWIAg2i
7d5y2diFdNOdnYNKV1Gz2d1kJYRlnGG2V7FmmRPwQO883d12W56Y82qTBexvqzuJbFhb37EZJm1f
8T6JqY58EPf8CuTCrcIhAlhg4ZZnrh3Hdu1UlsjgvtuM8gpaAiK7d+jA97Bgc+pk5BKGD9hDxKhE
ARza8FcGs4j5xEbomYAaQifJtmzMaGEYen6odHyjyq3b5dDBumqU9aR6eSk2/EmKaKAv2YHWZw8c
EBaRENq5nBZNn6C9PzI9Yz2xhrYawN3yhE6dpMe8Mp3bPo1mvHYehdoaNggDra9bC+XjQu+sJQEi
zDN8q4vZghY95xdQIerIksqcWrnq7HB7HOdp6HWIRvcH5ArioHxQbhnwZeVS+Y1mvR6MTbesRxc9
TpbbUkf1fBzyEqzkXaYATKH2Q5s8T9J5aBYeWOwtY43EDatRV6UeqZW82+flTym8Cb3VyWVD9Hll
5fVxekf1mW4lEj0NLY3Ql5t9gxt/kTzEDi69sp49Oc8CB4K/QV0NX8HJp7KYOQoVu0RireTPQZs3
UGgwy9nzwVSZuvE7DZ12jofr7dQm76uR6Csf7200XvTuTAydjGrK2TvwXK7CnHOursqLM952f8xG
moJZIEtD0NemJtNBSoywWMpuqg5+3RAUXfD7gwQ8nsyeo6V68rfnnmwqqrnSD7P1VRUhFdxFEAEJ
cBHaY4lM8gAsxdIp5hgIi0dW5bAKvQIwD32aRZfoz2x84iNnOa6oM1ho3Z6YlZTFGB+EjaZhzXet
5u1cRoIhTEJpIjgxDpxZYT+36v7zFnLLY+eDFJyM6Hq3thn4L7r9mAFXfdQ/xZiBTs0RXuT0eon/
Xx2ZWChknSQWA5Kp3TodbLrffX7xDzApcF71Qk4HC1gKQEfdeKbQP4WcftNQrqbxzOIYI2VYee36
7sCxJSIceztE9/s8ht4VLwRQAZ+WD7pFYo/mRH+L4Nd2+es0oLJFa9j3W1faGCVrXkH4Z+D0APH3
73G6tEDqY3lnpue/HHnWT8JjzzajpMT9n2zuP8WFKCftwjv5Fw2rGBMss0TluK5pRNFu/9jewKGR
jMogKCcTWY2B09uAj+7mGFnkgyXSE5hlsycchYbmzexymVxWgzpgm2ZK8MISPIrEGlqa7YOe/2XM
uccfp/yVXDdGeuGhgd01ixq8nlHhb8iRcJt5VFq3afx0b+rNiEx6Dbn/AaTS7xlcvJWkvU6zA30l
lMR8+REJVfmVjny4cD6LO4oqC23dAeCaXuJchpYUpful+AAd2bNakZIZnItAIxLHAsmy7rpenfGK
p3CFe60Pjigrf8uYvaCUqgdgzI3lxgqoEUSv0HjGUJSWURNWeswX+/I4aMUVucEGZVYM/a+3jEhA
wvblqWrZu+pIixAUWiyEePfGWYKYV01j/slYA9NWDYLQMg/TbmP9sKmnggX9K5upC4VLDqtLBE3R
u3RJdBiKCStSwpT8RbzYu/Nj26JznQCji5UVjuA+sp5FUcNmOxSVAm08cuXbq6Shh+YlcAoUMVwX
zGfsVWOaQoIeUtxCkE9CWd/EN+sOUUvjMGC+uYyBQGU05KeJ8T4g06aIPuVX+0AVFBGVvCwjK763
DYmY+Nrqinl3M5sPOfP9k1PHjPvJwyuZbinGCD3dMWlhTNFDndTtLwRLRgWV7VrFKDI4qNIItnvf
tIsyfkdaOxlidcVw2N6R9t2Ot80zOq0ZHf5rfmCw+E6B23VjDxhJFaRxkVgg5EPxI7qGU14f62Nm
0uKJyPPEK8dd8b8eUU9AUkPHPi8HaRt5rFfWLmQAmxTN8rtcJ3qJw2CgG/xGzPn2K5MzIXlBPY6H
ze1rW4n+F/38qe2+uB+VreaZrq98xzmg2Uj33fqQNCWZu0CadvH8yYiPMHKJqmkV8Mlp7WYuhsTk
RJ3YiEMAIyImqHKPX1+t/ZeR9i1he+7N/0wYc0opFVeAogZ6RQNeMk6ulvkRRXesvfenCl1J6j3a
X4sR3cI25LVhDUb2Qj2HPybhTZ3qSrAL0kCcOGbvX6a4Zq3vqLwiH0Gbph4tNTP2YpdVnAjmQTau
f4CdV9t3Ypp2v2MEm39TpDw7QWBGtxJ4HN/hHru52DSlJLTnDIOMb0t6CDKqCzf1ZbI3VkO53fM5
zuJw2LyLcwEI68/iidawVEUW76e+xICEZoKKQYafqDX5GR5OmCgI4EQ3TxhoHPpOHJKWa774BAmu
Ht53SwTgBr8hvnwGp2PIy+mrl7wnQa1gKNqxfA7EBqaZ2V9BDKRWEHNd3MTIKs0wnsSOjwg0SGf/
9wmLoJdxQnIwZZqE5JmD9BBlPgLjWEyIAhj0He5anJRn/ozo7+BoYb4hoNW8DGOnLCl2mx0mOc7Y
4X6W4fMpQ/mz2uqdm7ULbYzsXcTqmuTbraEh4DU4vv4T6Ss1dY/0kxK5sVvZMk0tGjE6pUvRJUYD
KMr4lKZ/AyLJAF3NQSp/1nOif2d2S3uNBB4dg27oa3zUE2uqL10ksFSj0rAOImlAgOQq3fPajmki
qTmTiKfS4dfEGXvaf2MLPThslceT3sfxOWyTVVC/6QZlYUV/7eNizTZuC3JMHlFsgxHm9QGnW7CC
3dmZAIW0oXiI7Te18vLfc9doLhCGGltcujEIfJyjjeiplmUazlAgTUloGZjXg7WJ4m1FY4ObOvD1
QPnQmQ/AYkPzippSfumUm1lw76A+rQIljMng+wSFrxYsSsNlnaMU7CvAwClpoeBsd1LaY3l1DoSQ
ps8aAYSEz8aLUn/qvxLgPN5EQR07+9D7KS2/6UEbhP5g0kX9DyuejXakBVta5cqP6UyW4+4Mzehi
oPnh1n99Vo5Q0NBl7X5WrBHkTPQ3jsefx9VPazhVnUlQ82wpNHe66ip6r4DkUwI8q8MKMg4HzWGP
a123Wiprnn9mbE4Eb143fbTa1vmwMj9111wr8VojM+qbyTbmxc8xPZRBBEYpqsUbfCkEOUZ/iuDA
axr69hcWI+2TtXoOmlGH3Ly/x3oIgMhLnDW3cMTj9n9HNlZzNS3Zw4nn6T98QI3VWhMFUj3ugUzw
91ZR+BrDLeCTpUvl9YQGCeLF3AHbBLk5luD5FynW4xATlDOpxx8b3bMGZ3OwdTewzlard57+YhpV
vUro9CIF5XaueMiIZeMgXKJYh4kNfPTNNOsbneG/KkqGWU5zfspE52yj0adA040DqWmsPhe0q1+/
VsOLvznimi9hU3nXeOttiIQgYWRifDcQWjBo11VO+RTFd393/kkF/9Sj25oWzfRG+VG+nn15eV+r
bf2py319azyVjGtMDZtQx2FAtkP+6PSz/k8cA5zj/X/mKjuEOx5H2wDc9cthjX3bRbszz7he5H0M
qNde4zVeOwlXOvpONJ2DHekU5tgSPXcY2PGs32R0wsuTfCly3Gkb676v/h5/0oi0TAIt7Mi4dDNp
HVWEtHhs44bHhmFPPqiAGq7WG/bMED+UvUUaA33emkXPzaUzrO1y6T/VwRvJsMetsy0gk8/2FFXk
/1MoxwEIcSU3slAu2VqAKgs9xfACVleQWRfeEgra22/xGjpGQ1sqbLjnSIUXDibpHeCJdYO5njOF
n10EzwFJLzMAnjh5ExR1qkyi5K+Z2H+hBAI4n4+UfYw7wu7jv0ivIiU4kB74OYmeRqTuydoYTheC
WH+qlnQTITrUhTc+/ZLsLcA/a8rVfoNekN+w+pIFOobzfMjGfz96bd+ONyHkQWNMpNUCGBfwYd81
RPuoGJjje8jqfhqpdgVEVQU8s1wGTmSFARoIwkhTKDjBkXyuDhMUoPTAG6XahpGr7eSy4nHMBhtz
jnNjs8lqbFRW7fky30hUbKjSMV9eZoXfTwfsqzv+PL9GrmH4NMqBA77HdCNs4GipFaPCbKlPfGu9
y7i48F8+vpjeMZa3FljfqDe325RzT3BN0cwQlvtMVwDt4tnNQeZom8EQFlsWA7bL+/kNW1L1e1m7
dKLuBE82d1ouAc96FzuhL+slVV4MmwGarYGMKAZilWrMhdpnpBS2hFm6sJA+OmLhGQQeFqHzLCxA
+9ZTqyjiNFw/po7dKnxW/yLtuUZkIhltGY8jfGMZyGUiQcwjc4ddHRtoe1bXBu+eTGzPJjNVL3Wq
hA9UphZSZrQO4qWyV8rLoNomVVeKtSYAvhi135A+xUlGr+abjoqoOWULvkOv0UlCxkN1olQz4Dtj
9g2YHHB018gWXei88EdNzZr0rQsMOjAfvnrN8MMFQb4GGO5QzdgLJ8wQUkgeNJjdd+TdV+BzVGVt
G4IR4qAGNi5Tr1X5w1Jtr1laQxLER5nh0PoirNLivWZQEcMWTlEN86WXHI71vEwW/BXzonjJpstX
WIYpzB0ZtlrdjSGOVxPhmECOZ4rMGX3znbCpdbUQ4Rvs2/Y0locvcRsXFOKYHeMNVagz7QRa0t3H
Cx95IwIdeoJxyEdI6Yu+rqe+vW8GWxJZIiP6f1X/wl/8lFphDuuALoMoGjfggrld1QA79o9OGSP+
shbPnDDtWlzSHCQJ3K7U7q6tXMzvc5QK2O1RrZ2A1XdtqsEBaLXaYxnXoHQmWdoDYq+A546Kh0Rw
iTBg4vofrNgJs7YozKJHi2TWrBj1cQJln6xTpe8Qmo3Na7uxvtACXo/qNPyCr/DQUTBbzv4xDzSD
gHkHkD/PWvEHdNxvA0PLVB9n1AF+hYtMRwS6O8xIvTc97LAsc9NWwaRGrLRmoXouVmtfCEE5VUI/
0TUdkq/pRv49Ve0Jmx0NVcyddfBcr0ByLtvDMTNEts0WRtk6svwDgoSvt8LVRzZDQcfSM6mYjhI6
985GO2KrvtzVCipkJUdrqyqGOxbB7ZgxgmKXgvoylGSmp6a7OtqI8QePJL1I8NKVImYm5shSwxoI
EnG0ATPbjR0nWnD6fRaweLTzIg/UFmg4JsPtdPiHRhd8Be7EyiQqbrKsh3oJknqyHzqf1VU2BngC
ICbI/1GlU1ulSrVg4yv83D90vyPpJDALDXcqdoJjXtsLNP27NUvlc2FsdJKkyW9v0rmkG6/oszLT
EyVIabVTkBU7fk+tgXUO4hpmS1PzYQWg3Ie8x4DL23NIiMvaDpXrlXMxO7FzsVMid0kIGhLCY9fh
hO7IfVEgUN7M6HDjMemNUKMSeMk4JU06syxJm36MybQwUhGYTHj742r/0+JiY3WoAxIuBWUpSCMF
pK73cqRYFMke/OL+B0hPMxgKOJYZvhoLKfF51tTkx7IEYruLy+ZU0aR4sAdvgBx756HBEmiG8lyI
g9Rmw2Jty+QLBa1zHY0a8Edr3tLcpdE0qfNPxaXc+ncvYosIg2TY/cguHI/k2ZtWwQeJCcqwplzC
dsWLGcCEizOchBXpHqmxx9bVWV/9X9kKO5LYmiY4xDattgQyDgK+hEZD0Szj8HJiVQ+X/2qq0Yyh
hsKL75wAOCvueZRbfKIzBf7kedjyU/1lJj34ztSiIzTNgv9ix/TKcOjFsAKzxGspLnSpfWp+iAH5
2rBtlIp0RhKoWl/KVDMnyTiuo8epg6KNc4HAmRwYbNt+RCh0b4YS9FSyVtjeWvHqIqLOdwbFx2lc
g1+n/2gJezuOqS57tUZkCT/VwpcUbExGM60apfiVeTZkVzQt2anjlVx2y7XvLDj7K+a0GSFVW2h3
6s88zvQDIsaNIlK/t+3bhktuIypgRkgC58RkG7nKbTTHO+AJ41zxBRDpuyWk0dR/cV2u+B8Rjq/r
wDqtlYHjpoXQFSHYHFtW08xQ8IDvc3BSrymT7wRCb7BwfgHxKhHAvEua71JeeluWEkcou0f5kna5
3xMbEWdbsrGhnc3RbxdMa0hMkgJEeejJj4dZRjw4zm/6DzVCFSbdRsG9wJ4+XU0B3izYHtEUzoxR
7dSqS1P9gUz3pURJPOeGtscKbMRMhVxhAuoVpu46GSufoR6abpkiq2tpaFq7GQoLWngomm0hqifN
eCjE/wPqaBAObNJ/JLnSEyheeHeeU8a7dnFJvHgw/D5Vb5te6HnZdJSOH72EepDRabtLsDzjPJZ4
NC6QRHtFW+b3ATaVsuB1Fta9STrCBIFxELhuIrPiYKZVNozIt2yidMwJSjS8/FiExEA3YoMWzrKy
vneXIoc7A6sVdDgR+baXzvsOuxbKelswdhKGhIfRwm6IyIkSkYUMpezsf+YHEjhImroFEeML+gET
ME/vvwHJFhLWGdg3f5nuJaTu2A2h0jNW2h4DQas8JYs/x5NKO5AE2QuchhIWps+IxKWhwseK1qPZ
RjLu7w+XpNMr4onEUDxkgjE/D+B5575+ZJByQXwCvoTKaUSqteJBpv0EtLAhAygscks4Fr+s4prr
iOrOYcx0pdG1bkaYfAa1wOFbHK2blhschHd/UMNSflYXCTEfZOzsUTjlrqdfGyIwetzrmuS6zGvE
87pCbDu7ICfkF7dw+MJMdGtJ/HE7wuBNbNyvMujy3wfYIg/vtIw6nvYP/2pg9zBfqH8QEGUXlqux
LX6xzLvJAbVmOBLmhvkELnzWpAdMpd+srIt723wM/jTOOojosypH/LC42/L25eAD3A0oO/cz2dcg
h1xn32P7XuizEBtR4n0r8xXvwvczqa8Kqoxa1vc4oeDfiAih4I0fDmqyW+GQkuT2Uel8DKErZM4h
r5rM0c149HWrJQNJutA2rQ3+cgS4XST6jlcY0EXgIBkvU2hTNFzX9hmYgn2NS6zxkuXbuYryJlHS
2eaF4hfIdvKqTswD/aCpsKxy2VIySH2e78gGU1DLysjP6sZZ5ayJNG6cq4nvVS+bNggEJ4czjp3+
UrrY+JvFw0O+xhBjVPae6TwHEKvWvkkNx8ztbQd0O5P663b4kMoPdWZBW3CjPMxdEVnqFmOkvqhR
7cd9jnLuoPP1yHOP5OKpV4lbdudqqs7qMgIQiA0MQJDvEsmQO8n10lvp+NkjJqiXAnB7j2ZcCR+K
TfjFrxL4hG2KlWsKYEOyggtNBCoK4F3qfogB9l6dOmwpKvrGkbznfwkQg4zAUwRII2mZ5fidxCwJ
sVM+LuI6mIeOQVQLknc4ba9ZjTgAGdlCkXirurhVnfTFZ9dj9KChkIaFDfYRMALb+qu2cIkco2ln
rPEGeVEQWH6FuoQc7Fxmz39vnPahPqLVWYJ1wYLsLMidqIvQmzU3eOFvULjxePd/EC/0ozfWvL4o
UbfUWQS5OxMjcRDwwgg1szaIeTwoVsTRrrWkKUSBV9dHlCd073vHLphVlgqFeWSbbjn8hu4pHnQt
QFB7VWSrsiimkWnhmerrsuvSDlpVqna0x0Cc3dEmoWfbVviPrJeyOCnADUSheLS2G1pafbKVUnGZ
ihFQAGMkqZ41q//J/CQgD2uWqKNKLgtOtJb86VH9+vIiOilLdF6Hygcg/9UuOYdG5xArjb2OPY8C
tnkBX87vl+g/V61AcltXrpvXDLs4MpX/9r7JFRfCW+I1m+6pf3IVbfZ/FJBLJLFFSA+5gyEIw54g
JXmyNAMp/5ZaJQ5t1v41Pe16P8dWSVzRCSWbdr1fmkL8wdFMyCvqtubIil+twBhBv8HdMFneBz2b
XC6YCmJA4YuqbgjURw4f14C0um5h9PuHa7sfP3j9EhWfopqFRIM8+I1Whhl80k0z0oF/RgD6JhJ8
o/Wdf8Zmk2KqrX5/DBq7tmojS6WmH9cDeAXq3a5UmSr3ZI1O0zs/Mkklfn9jDfiDzLB00IOOHXZe
SUnBnpIbNCc0agyFuZWZmnzX4JYW2W86hGaDS7gyetT/O1N4dgZ4ewRMUQGG5BJpDYPHtFeCGliI
rQfUNBwBhLqEExTCzv9cHrboOz3CTQepEhjf6DETmL/bo4y3ynwSlnQzrQHVTTGlM6nEPWJhqLKg
L8UIFmQZopZozsRGA2lq+e5IGr8NKYtSi2dCf7Hsd6yMCNr2PFOJbSfjHl5JZdcGnseILoATvfFU
aXknoGZEgvuTBL1QJJ2lAm8+6Mkrdzis3Uu3BG1l8xdS7Prd0wUDnaP/RmrtBB1vKg8TIKkrElOO
nLOFHSat7APuKUmb7Y5U2DzNWmBV67M0aSr7HpdAUpPe7OrGFwlJ0X4u3IUVBG9JaO58YZdItjZD
H1M0lPevCuS1rwFZ7z4fcyTwfx9nv7EYFNqys3G0Y4+RFg9XqNqqudaxCEAQbTNx1nYlK/RaJdLD
AP7B9Rk/6Y34yapXEr3HlIHHw8loKGTbodjCn6t6nXG9Zegakyc2lfdm++08M0m3SUFT8NR+N2p7
dH3yovzbcVmyXWMSk58/kk954l46ClOHbvYKO1QB0iFaSefUOqQ9AMq5WmXcKxy5Kxf+NaST+p55
3PMqSYyHBzEcAKv5qaSfgZznrQk1u6jSzfw38BRz4w+jVGR9Y+7AveXmLKatbCSjHN/3skoUmAJ5
AeOYuAPrHRIdxUwOq9xkkigNWG4P7+TeMIfPiyjMlwidvlJ+TKF69pXa1X1v+Y4TwohBexedqO1O
F5gGeb+F60oH8NC5I8tShXnSH5MUrSrxXYwXb3J6SV02aqsZNHhSD9lvzLJdkz+8GiX3II1pSLYJ
Ht5V4HlkfxxFazakx9RQnjXXcumswMyD/qMPFPjCHe4HEwg4JwUUgtWMr/qlj6w/wAuLkO7s1BVu
FGh1RTesA1mrKi1efy0wHZBHaF3VbSK8Re37x1iVcNz7q+B1vMeal561M8OZ7DQKaA+3qFArDZnU
j3Eens9naY9BP347ndl4woG9hvW+7dD4yjNd0LFLsCbVWNjZyeEjKMMe9+50jyjC+n2HLLm2pY90
tc0ezlAO88azUuCgZ0W3mbqN2+tGNvOy5IuBjpPviOPc/G7qcHw1YsL54f0+KaIdOxg9AHUBtvpT
8O+nXii4e7aV+1ukKIme3c2cCMW1Ml/J0HPI8H5YOlFOBCZ1R6iNOp71hvXaNPFs3He4+yHsjYKu
yDvGxrmpl+bdXncva5TDh7jHRpzT7m1L8Oxn1x3EnbEqVzFPM/mwGiZemfiUtMQB+t7mhqmc4jjM
NICoxT/nvN6+dSMRLS2Yqij3rniOhW5CEaHseJAdwwpOCH7QTP7jEzziYvuaX6EhjXAoIh92kI3Y
Y4KbaeT3J10ygb9cwjZ+aq/vLRehuIbRb07sCAwLdJqGNPM46qRmOaFVanlJGrsQk3iu6Hwj7HoX
vPUnqGNAIUIfgCFe4XQ9MhxNLiCf31BMlniEQ1QSLq68nEUlNkIz0YetkYc9pcSbDV3KPYwQpxxU
VG6bpES/ZmSXsvHxKLsMgExHJpEyQNhRxUjwb1LpfGCqrncSNCQ0zWLkRBq26RkzQEvYk0b/FlYB
XqVzsx7YU2WCoHjK8RmTLZo/+aLI7EOtU7JAkhCsqZpdoK0cHMFGzoqEZRlcpRowgJeTNdSyDpLk
m5rbJkyC3HakGhyIBzdwCbGoIrBpRyNmj21MnWtPLsYDiuw+jKK5q3JH2hHUdYEmklT8i3/Zlxsw
3oseaMl+sCdB0Tzdj7HWwTxbZPzXd5yIR/WtkBIQdXVv8RPxoSzvA1x/WeX8O2ohsI0omkRW/Ogh
RujujytwTnENKUcZLtgCgol8qknSsw8V2peMAJVWjRpUic256W36sgRKm89DL/3y1kaX1jv/o3zz
FBJC3+kXosP5aAqrTYIM0GOJMBUl3GazEEIzkXOymVouK8hJyg7pA0+955sCIBKdrf/RL5koJ8P8
bhBqKpsS6f0rKmyKfjysn4KlfSKIc7UwSBeywrx2oIGESn5ZZA+jGp8ER3R/zbhaEdoOZQRijGCG
cGozhwtKVHavMSL+v9prdU99CIK4vPjwx11wmholasK7mjYkkDTbnHfUqqeLSYAXAboda9zM8R5x
U55vSVNYSWCh9Wi3jHTQPqLDvuvofCIYuLyAs40FdI4Dl7G7fbfRnRega/1qPS6vHd4fbfouXRYl
38u29Qhz7NZzSHwrADpEVXjfQ3XlS9bP8E5Q5DYH+lpnkDtlD9Q4UIihUZ7L4tMAQq3KVlpZUQbw
G7ft9EDcEzeaXAVFGhMS0xyFb2JsqiKxwecmVP51B8G54+jOOOFGZvpj8QVWvjACVTVzk3Sb00qX
is8M6UJu8BA41LjMaqjIs6jrDfyqwJmOATdBN+Dw1em/PqIihQoA5KH7XJbl7XVpk9R5X+7b//Z5
CU6Fft1oDRTqcngXdRREd/P1QIr6aJcJJvNt41Ci68EsMaBw5cuINaVqdNl1XbD3zCYOvrmNYdnO
aMlNaP0amHZB9OnJRtfALLn5qtMjoaABOdoiYb44wbhidEsT8VevqNQ3ARDEo8PAUQ/KJ8pvseh+
zUFEwalAsXPHsdipsl9PkDC4bYcy7nmNDos+YBI9746ih6Y+HWgUgFldGHbEhCh/HIE2DmjOf7BR
z2EjUFMzLGzAbQi6biRucx33UuedNY7oo2UTg9xhpzZAQMfYDIWaSBtX3fRfgGGoZkjvJm6Rn72Z
++Br0YUEI0LPRwb48iLy+CXa6vCRg50JcICT4dMp5HKzMcr50ZUiYQvK+96/TIZuVfg780YJvcKU
3b9yibeuXy397EIGmZ+C819TjmUlX6Mo6nX7ERK22cMM6XR1cySMreJhZ2+1fC5nrrl1CNoEcVn+
42jX4WqtMzvtZV/BuwR7WoBVuElarvqLmO+KuPSFbYwBkppbWK3YRBosMw1OMNes38LHYPoZ/mIR
oPhEvr4nAaYsh2cdedab7PQ0rggR/hl1PyFZVvgRzzDzRYi4diKxHYxkwz6ModmpARI+aci76biz
LuWxpq+4OPfcrSY1IjcTghphFNBf12/0ZP7nt1whUKROZ17T3IpLfz5/wvd+s4yLne3EwIz58qqD
b5CQ2XUEJvZufGLvGkm7domOkOnTFi/mHQaCFggb6uqCqCQuT2W3v/Kif6YWzo2sWdgfhvulX1+Y
QPNMCdXKv154+N69RfsWVz1dGw/FCuxXAWxztgCNPi0K+VBmTj/Xmmf/WOZahh3yoWyqCWn1spw2
e3cA/8eHb1jDBQq1oqQCo2eF6bn+1h9Ay2FzsvXtEjAvUPpi1p1ZUdQhQ3B6zYXa/ZMzVpr9kwuj
6EQAh+u/XfHu0LKTemIHUD8NBQKmDYHBz9XLZiv6F1VR9g0maEOrf/40sHGnZNwn9R6gO/OGkZ28
a1H454PbOEjMUkrwokChrNCnsq1q6YXIg2tLxiII/1ANlEJkR9rnAIuoKImc0ZTOtKLUtlhppEW2
9QhyPiWB2miKuTDrDGPMHSIhz/Sb+aQr2YcMM+jGZChNb5Bl6IdjfOaYjFL7AlTi7lUW3s7rN/qr
K4ZUx8/5119CS4hsPGHig0X1Kj6QF2yP+2JDBnBhUQnEulmUimhi4e5GU0zodb0mJATOz2Gg0FJ5
sx0KxAfgI6vL0TG6bGJE3eq7Ia7dBCK4In+fI/5W6IjhJUozR6oHErj/ZyQKnk095nAB0Ut9nvME
iD5IK5Vaa02taS9lOgPzaiikmYAFe9udmqM3VNiludpKnve9xxLJlMhexfdrlU1sYKJhXFxRlztX
FVwGjo9h+oHnq/rilnDVz2/35F+gDjvKB/JluvmoFJ7CIK14+4kAn3DKLPZIA9AKJ7TRUSJYvSmR
RxWnt1H0l/1qNoNAcb2O0nzlYn2CvzYYcNS73rDH2n4Ej5lt8x4ckwMRDGkeYn8LQDquJgvcNkEV
MJ7cOe25cg2git/0Zxui5cfgaINLKz4pjcWPQO122ohjqxglhZJHZuaUovd3txwNXFGtFBeQseI1
1RaNs0LBfMIegus9DBjT8NQSLVyfDGOy1bahkyy++UEdP2e54Pqs8c7QjUnQv4hnigWGGR6nJipx
maqr8WtYz6GoWWw6dHHDAV19MOCuIndzZvY3VCv2Bs5qaaqWZFHCD12hQ0e4KQ80mbafKW+ggo0J
2FlTDyr+1YbFM9G5ogyyoW6SQioU9qy4pE81OkYAQiJrKb7I8n4goIbukkWtaN3JHwO1L3URO3hK
MnC5YDUVJnwCYpz2NgKZSq1L2fJ5wskiJRJEA3d9JvEm9LvTVTr9yTZh3c7RvcLyLT0p9wFvGWWX
bm8awm1cJ4RrksOwxZVhBaKQTFRmgXKd8x/Kh1gO99z7a4S3Cdj0CL18brbxTBSYT+B8cc5NrXHY
zncfdNXaWPCjQUJm1w0aZ4QeSfPDuy5UNALjat65CKq/PLkxeJ5VZpteZRc7kdHLomqvmYfWSAz3
dUvw0fmF5Dy4o4Fr4J6eoZ/0IXo+C5H2hnMbI060ArzLtbUOUyebZuLn1nRjOLh+goniCDHUhi9c
tMmX6nkHINqqn4Ewv3ePN019I4OwiAR2hq6pz3dJ7nAyJwnWOpkAzVDFre125ZoJZ7enJ+FRgXGI
kPztVkA22bBgImeQpZ1rfPHeCUWo1t5tnEGTbeseFOPNXj+HTFGppzlQulJmShtKLmg1HHxM2yvD
e6nqPgvt8oM88coD8ifn00mWFTaAZrreRQA/uA9i2zwtN38cY4nC6Kb1COaeKtwhpH1qxlLvkpBF
AilAvPONF9H8k1cBLZmNFZR339gh/yBllTV7Mw+kObjmc0HZn/HtmVeX2RimPBIJmIvPlLyDGgE9
uxdAGAHk+LxvuH3QgxHDSXQ2yyA5O7f8ggfMYh++ZKNgBDtemXr7belqhuWP0bFE2wQG+JFdrj/P
pEYVvfDHfRjGutcHgEEISIn3KFam5dteRkTs3RdrmG4QLEvD2ie9+wS7NkRXc8XyRrvmXLt8jWRL
zAtEPUx8cY6q0r279/ik8yUmxjn5Q/+z7fxlOT6ShNYVYcunAr8KDpGTZg03+ohPsHdoLiWtV55Z
272HKgyEluLf0kO1Y+sKUR9XcJDjwlgWfHOrfkofXTNIoNxrdzfxmrpa3EOpMN2ZWG8mWMhtyyWw
sZ85Odnet+Ec1vtesUN4aykNW93KHAIm5pIr/4uBs07Vwj5WTECysRPhs9XaFvrHcUPpSXyXGFFy
DnmPkyBPHR/cHY3b1BIFDO60FiLBT3yxLFext4PJuZRun7Q+hpLbEwMQwbXxEHbbRlumlMAWFpzJ
6Jqh1yG3CfVw4MqTdQ9e7S2SDD/wx7RVKukMitiViP3X7u6lX46Lq7418crmL/wco+9opeCOa5AL
k5k8P/wWTs72c8PEDfagFTWfAg1vQkeZr7zo/hEYjeKDXVbRbSPlb/gBiv//DHhOAtphFkMjJOMm
ImVwKLireyll/Ebp3dO3W4Gk2OiCsdMHBvuuD1YqTMA7yRWbnzeeYlwraQbhi2ra9VqR6nfEJUzf
WhNG23E42XSkzP22LbbNWqLa3RffPNmAZbzemlB+A2L9Sry9BomaLi88K7jYSq9v02U3f7r7Vph3
h5U4p6uCALusJVtVVJzz9g4mIu407HPazd2p+TuGYtB6OK9Yojs/87uX/NHhl6WqIWwLnnH7hToZ
sZbdk0HlEU4zTyhzX2ZvtffjF1FVTGfAzDk8lPl3zOCrp8msRWPo6Hrs5pPZRKqXMD9lpE6GX+y0
YKDyYGsJm4WQzsEReKGaFkk1IvOqvnMVs4OPBXRRQio23J4GPCO5EcPrQPGK5npa7FZ6/jA6VjA6
gb8WNSZdCRPR5u1imOvQLmmHH5LaO9/VLoPs0EmQYUttJmpTgBVyIUe/81x4r1bc7VgSQid78VUa
8w1Ii0FijxldZItTH9zrglM6JHBYdZ5T8u3/s5OdWy3jJDgLCm4lIVBJCmtb41HAdloFJV2wm5z+
t+7UwNzlNXoF2m/oi3oJxGK19BWqBLxOZhnt2lqArtvxG4AMulbOHEBeYsrRBc0aIGcpO8vVx24N
DJaErV/L9GalSZoV0WXdFmmUCmBT2Hb/ao1nJ95Gs3loxjxLWmTkP9SPuvHWCGJJXS5cadVQwX6J
EgjCq7lYKXNHBeHbg7XuoORc7yBl+5cVoPW0ObeYyspWzYxPjG4bTXpKfEabAKQH3A3ScqZYzYLs
FxUcqOd+YZLbm9E+q2YZhukn2lcxWvtxfR91Z+CWBAKXySiW7AOW6IV3uYXpUQj/i7DM99PrFKcb
kC1m8JV/wpTw/VeUP3ed2STjzg4ooCrFxvfffG4LyB7pe6papau3cTXT2DlKJLobouvN+RSsHZZp
J7PGvaZthSxFRxnnS0jfsBMUsE1tcYuUCImWMdEcWUahOOoGq0gvYkjdDx0BPDVamGj9x9SmoOcy
Bxx4lHmzSE7UhNwwTTS32NgRl0Isu1TguRUzEPzEu5ao3K+9Vw1DgxWKAzfF1uO+UZQZ1SSEbXCn
+YvAaSEod4AaJk+Sch6ZBx7KcmywhYhc6g+C2EeYlK7k65OASw0CpD5kLFGNYitUUTvWotFAQ5WP
BBh3WaxvNZUuNtxQ5OddgMR19hzZV5LI8Ky//82M14cLAyte7QcsFix3DHP/xeUkl0NRITE3UNhZ
Md1iqpzTuPZhqVWfIAEtYQsWL3ywEpMjjnagmLWOln6NkEdl1+0zrTwqC1iTPb/R3yW1VTPNw+To
BPDS6qLk973x93xp9TdcB7Zp9bAcIQ3tldjiRbgK7o/ql8Z0MAVhC5jAf3iKKA1omS9GM0xGXOnA
oQy5iXy3I0k5xRu42pN1v2xvcStHiSIequxDqQN5Bjx49CeMBgRg9+rsJWlnR/NNAjcgFgfgk6SR
F0E58NlC3+fIuTF/zlVhyK2Gr39rhCj4fQ4KNHGQgMrAKXAJDLQqcf1WWLc83tU0zS7FMUEhhZoC
O6Ig+MwKjCz78t/Sq4+U8mnKOOjJscbbC66+Y9QOHR80z2fOJZURmMVZ2dIb/m+jojT1K3/OAy7B
h0nBV8J1djJidJ+0cxSg6dpOQrkN3/YMew94mqyKxoG5F3/RZCRZDcjbWlQbeaf2sl5PX9EINSOs
90fKmgWDha5JgNKkJZCZl7MQh7L+hMF2tp/AuWEi6Do8NMYrnj8WnhciXVjfIM5AX4yHIBuoZD7c
9fDJtnWOzxsIE1Tfhis9O7Gy65CKthSqzO+ksUxr69weh7chRvvMpLPElJt7W6ZE4dZdFmSNV74/
aWl8BHbtATzqM8OKTlmD0KmrDM5G5BxT2Eo5cZu8ftPOWEyTyYL/pF3erewUntWj0088AfaEptYL
AZeI96iCI7kBqSa6xqF+uEjkaZqpW5dZ1w8DENugdjPeoBbyWCTNl3GYMHT6UnIVs2alTMOnLdPh
fS0A2PRlPAz4qj3IFyU+BqviQEvH5jrnFqCPcKRwGehNu3boAEPY9HU0WKkXtp7HRDF+VlhU8FUY
m7ZBZVCJN8I4Q0Ddo/deoRnYZ1J2cT+pgxukos03OSyatO5oF9lvpwMOshkL47MbmmyJkVGqhqgC
w5eiQ2+Lv9AWvfxSdbfFSk760rglk6Ut4dtcEj4rNPTKSkO9YVGtbKxURw1FlwKuzvD9SOye3NCZ
+gGkm3jz0dEghS024XTaf3LGRsS6hJjXNUER5CH/HS/vH9UUezPeJyxpw61B73A0m3A3OvtEJpUL
JZYakHo4+F2bKLP5l26uvzgDhDCJGjtUpiq0U5OUNv9GLtU17MgPNiM8AHjS/GBMS6tpuz8Js7lp
u0fhak0ylNVa7zWGvWrH0kLzzfpB9INHP/75F0O/ASaBHJCjS48mojQ6EwpjUhm90Cai14ksSAx/
Is81rZgij8Ao9hR/QHLV6yB0+EZo72nt4OGcKf9+AMoxcjWbJDbAyseYPAWQdAvvA+gVeUwHMHyF
tLcvGeSJXMYvaut76J3Ja1mdVeFQasbnnVzb3Jynl8MDOJlhnqcGCx5tev/81ilCsJrm7wqDaZ47
jyHELxgyQgSa3iBGdnO1J5mYy4JNkOpIFSaRKOv6bR8fwQrGOn9FDlN+Gq/nNeSneAcAYgT8TweL
Y64/aTYy70q3z1ggvenEj3GtU7Z1oQy8NPhppEaDWdBMUAWy03vfWaEouJ+ry+URjj5sBVmIV14H
G2xjSpRbkY2Mz+683dp9+S1u9j5LlppVdLgI3ZSGnoTuvHhYQCE3MSU+4V0U+W+ScCiXEuw+BZca
BhAGOydwyb/YlnX6EqRW/SwLJsKFUATpQPUXuWBZYg6obok5dj5bojuluPho79znS5LC8vI1fbmg
9JToOWDokAW9yjGR4JnLQgKPHGRAj5pR8f0Bd7p4By0ZatrXq5m2a/1nn7ljV43QPd4yAWrr35m4
20AGdoi31OOBJCjPf+CDn2IHnWiHITRM4RD2GDZ5oeLJOj84Jw1SaSAwWH0nx7kxcOyWOyPLJ5ys
FUIXiTEpSSOyS6MsTRQnARBQYupS7ZDcUF3Q8mZtPMt0KLqFkwxW267N7HwsCBflKr2qsNt3zxo9
eKCWIPR49wJEbOZXTGMu9OHXf2dqxHTW+TfAzzzkaBLPL13iVmQiFzoKbRrvYgRRCA6QJp6tIDVn
EujRQscfuuhvHSPcZ9eYw02P+RUa15LUEQXKGLwfFSnsT4AiKAAwqfmPCd2zxScUMV+cM+uYD2Sh
CDCA4Cl6BdVyfumQqGvuRKYlK2m8OSnMEuZI+K8M53LlkRbCxKyWRzKgsYbDATyNr8MWMZR8TJDh
PMGNxPRpTs5rzoSZ8jrmRmBynrhu/nm/eUFVtBYm/6q28BI51tdQcPmMBgM9nZ1U8svzlgJLbJLR
D5nLqt69XC5mcCpQMcVq7KWxgIhPs4IWCVHuP4ubrAzeqMsG73xPtQnOFeW5M/kMXK+uJNs50vMi
G1VirTFzBpmyat3CuPA7TwGzX7T/yx3AS5+fsKsB/tRB1wWwqp6mMMGGn3YC9FTk1g9Ydt49YzCn
YqNdKfFJNQHSxZJaO/jv3z8ipVQwUiMJrfORE91SgFMQKls+3GCHrEXmFYmVZv/fQFRh/8CrazNi
lCea4dFQEbZRV0T6a+4W5hcIFPHt6eNQWxyWKuEKJ+GM8k70dEGDRKVj5IBqyZMIXucHBhdrZJBj
L1iXJT9+Fvrzs6aVMuO2go9835LnNI29MPykxc9n0uiJGVt+FPTi8f0aoMcT0Yn2QaFNLrSeV3/B
3byykqE6I+YKFRYaL2gPgIUbbw8u8H06oqbIQJm91p0dRAb6LPp7oalddN/LHHqHWs2EtGxEzb3+
RJnhS9SkK1Ei3JKIGs6LoK385Xn5pafMc5Db49pExkLiQYUWRByKy3yNHZAGv+pHLVAnYB8J18/b
/UzTCUaKggrILQvNhnBgJPAoQzFQrcCAscU2zmVgfvtALbqiLU0Ng5rjgK4BdYMJpA1Oc55UVzzn
5YunLWzOe7Iq12ppNo8YILxsiBgDkvfN/bJkB5TAeDPsvx0OsxFbJ9OpNbb7+8GgULGAfZFsI3U4
9noissHYl9Po2vMAllZ4yrxiSiEaIEoos3iqi6TXCwo6Q092Nkz6gwGWTgdSjD13WwsKWQi/L69B
NIXSt6FV1qIc2WrZGAvSzxJkagCX4u+x7HKbe+/EWmIa1+M9LDWMUsxv2pE/058J+2M/lxknK+fA
UEvVvDzXNPMhNxfO2GXLU6TPgIldq+MYcT+F0+4M202LD0/B0cy5uVvT4PNvHx6JeW1Homr4qf+8
TsR+Z4dvLRvw8OxsTmGwFPRJQUeJ6KYwea93srP7D9S2rVuzDiMh6UZirtrXK/I3GXnBmzkDN/tt
1ZJ+vIy8MsvYhzHJtlPfYPwuv4GKjh8fKNqVeYnt9Tjdgtu/sXzi3QPYm/dBcAwCCGG61uhGC17z
y/XFYK5Qd1pwyOMPBQPsgTQa7CZ8L1JVZhz4JJVTNuKHGHXRSPGlFoYmhbjunEzcV9GFPrkcIyfC
AjtQYSN7BClFRBowLJqmWkHXtFrmn8eLtc+xp1Pl/vuFtaubWY7dH/67OFefS9ypmiY6veTzV4K7
XUhvfqscPDa1p6Pk53Ir36J5BVV5Ve4JasudbAnvMC2L0TJZynoM/wjoDj3F9rDaX5yInyu3/kwS
+ZxzvR3xh2bF9RzmD40AYtdGu8t2lNNEtADimvfxn4wDZknnJMiSr7at//+xkYJ1BJaurxae+Y4R
+UTv7nqrmzusBJ6P/Ph8RYiQOqKvNwt0kwMq+Sl2kGw+kh6V0etiyQ/LAFsb0sDciCvmQ/hVFUlm
O+17V2mzzjI1/n7Z+5jSTaCfMnF0M1GghvdZMNJq6ZHMF4K80I04mKBtLspwh/k0jlA+W9q8oemb
jrDdeODfYjXsk1lryRE85aD3mvQl0Sb0W7EFVeoCYkjQpUcJHsRdZw1RTZ+f6DjbFMKcqRZHqTNl
f6ogDOrHiP18qeWSyCEi975HOwMaImvbNa9ljpTNV30nZsd+UxfnFbJvN1XumezT3mKnMEQmmb6+
QAj60qzPXhpoeFkJgtH5XQhfMniMDYgciTOB7a3kWdnAAAnNW4PG4s8PEhEBMAT8EpX/F2QaL/bf
YZOeQHs6D2iFusL4SUsF8TPX4oNyx1tcwPNLrejP4lao8SNxNVGXi8TN1txiSCOWoAfAbGIwe7L3
CgW41xcfa1xgZ7+siM12YICfAIwr4X27RnJQbd1TbGe/y4IuvNTpkvFOyoIyJflOSnEsVGkbitCW
ImL+jV34Q67ilvzmhajc2ZLemo4gsVgzWxLoY84aiC0lVwcDASSeG8DZs09T36x9mjsGYC3T5grP
kdf/kI2KSERYGeVuFnpaIxnGxDYdwDZS/iJof15G21zRz2U/Np1JponnE99mwJKtBFOZyJh/gevW
ZUJSMqJOJ9/eiVepEAjw88ntAQykyAF1feVXqa0oYwcCTnTOEEISUOd8WQ3kedcy+t/q8XungOQj
kuR97UGbfB+2Q2UiDyEKLTuN8aBxOVk490OjTIhtNlKe49OG8234E8QJ7SARq13STlQGDeULUOvI
CpOGr5NDopvxXTu1ZBBY1/25T5qiHAcMxdvFzfiZ7vvAWt0IHiHIaUt92R/esRalM80WWVykEHR5
nJAJBkoRUadqs1C/mAwVhrWS0Z3LeQSe+sMi3zJydJjbdf23i5mZBJ6+9ZBjADRd12UrBEDKW7nf
sR/K6YuC4Lxtm+ekBYbBQUtmawM6YFPuWeRIiZvGenPM88vXWbsD0pJ3HrxYY4hsPvTDEqx0Yg7R
CiMU9TBrkpcsctIGosRUtZXLhPgPn9UYSyVcQjdbjWExATAOeJTc+sT+bjT/m1oMj9P78fLJcyhR
XHpcARJ+a1/K+6muvpDTPfLCLvvoFrWMUjzjU799UDJaHK2Zb5F40fM3uIHFYgRjpi5uON2WfRaY
bQVyLE18cAmSFPjH83J9x+Hy9Am02AfLgXC47XBh5VV3tD1VqdFuVIGw19n9FjBCf0ipemzVL/o0
xMZ3af1St3r81oAx25szgl3qkDtKCcsT2IpdeaeRW6nvwNJ09mnX3z4Pv0/CGbtBV8pmFy30VfVF
xhAgtcH36uRYSwdFD27hjMvg4gi1o0w8poFIMeOp0Dc6p6cbEN/FOn+kQDxti+ymCWPkR6OQU51z
v+Sv8PxVnTzRcjD00m7w6SDEzDdQZq1zrZA52ymsOszjQLDRK30uC3mBk1OK4Z7KQyK5y+XpHYQ4
9MW9QwOfMz2E/MfzAJs1cSPhfrujkzMFJvGoDANmPlzkIlouUfvZgafNk+ppQw5TosrmO0VLTTTd
XvZc3QeX2/DifhWuptYwj6oGaJqX6DcMzeonuUB3yLaqzb9aKXXkAf2mggm5SCkxHxiwlFlzCYHr
Vf5f1gpHio6bGR5jwbTJ1Kb50EAvYVL6U0Il1kCudBIE/ucGmO0jqHqj59+Mkgve7AmeBPRVb7z7
CT+/7X5s75PIJNxWMjFeSeIbVoGETU8pQUDDZ/GB22LhZMB/zD5pBp2Pc4kV3UTk3+HddRCmWFl2
9tHf9jnb+5UIADweWcOH1G7mFP6jvz87ABSaXolyelnFI5S1b9Q42Ms+joP1gzv4hbdUE2b0xi3E
eVRmAm8eR4s88/WEHnJwGiZe6MW04xRytF7jRZakb7qZvjGjhYK/IkxNn/Z3SE4vt6SU5B/K3tsd
kQFsXbJJxV7SCVfCwujGpZS/R33pzdcFUkpJa4laLRAF1O8RFNDqEPNf+0wZoFxMR6ueXYtG8Kdn
8pw6VV3+kcK7NFZSAVchWxwQcRZdrWZ7ApZH8iXUmNnA1krjCEf6pJRVBfsGDunYE5WvtHMxLtAH
9TlQN0tDrMh8QfOQME9A/RccRk1f2PPqgA2OvxHeHkRUTGmtQ53n2Na9k4GfwH5o5nJu1jvwIw7E
kpWTRjuMUN+0/k8rVeBefiQzf6EGj9Dgb/ZXlrFUMfSQ83G0qgc1EO0e7eeP7GM+yv36niF5TegN
eSPAGZ2Y+umUz94hq9+bRiAWyuevoLVgVF5DryAJ4i4rk3A9ZE6RcTfUslrTWlYUUB6LMjV+4wLT
AFQOMZOic6Xu4NbnkQeUSHcP4DkSFviR72Oar7wQI1mLe11FstxNm2OuFtftWhrYCzo/eNcnRoke
hR67XmDNSEp7oQtDKt/XCn862JIqwx43NPmoW18/u92Gk6ZH0TWDG89kvt6Js1oBSXYIc8BXw6tS
XtuDgeHjvc3NqEBPm21h/vTTptgomLF2YeLhEdqBf4BDc/IHgdLs6z4MLhwb0cgIVqkKr9ZrvHOF
pPIUoDiFPvSVk3OJBVaI98BZqYTm0DHdoe7mtnkKYJMLfWwcx1+BS45v/+vfDNwcUqayf3R845jF
zofwQRCFKgGUH8zflP10kgCiK/Ah4QObkKRv3GErzWZQa2H9PJosG3RAz1PdtAwUOLSPejt5MG+P
CCjMMqu9vO3bWYzhaEeASsCly/DV1QRbAbBNnAZnkb0+UHDLmzWw1axSGU9smX8x5IAkCxh4AkDH
m4wmUPpQGEw36JCAqLdTlHg2Cs7iOdGXI+/8SzNTYyZx9l9NNG9mvd294aRLYDAGGzUZAMkroBpP
vmMQvkmboGpq+JLDFi9rGeZWjKZC4AVtbZzfc0FfK5/KtPi9CqhbY6+wD4cSTaOfZeWJwjO8O8T9
5U3TjYHzWdvEUaDgAZ33M052A5GvO+ztKMpW10ka2TyupDHAr7sDIi4sCpObnXHjWch3M4PNGeQ2
mBNX8x4url+uqHAsul4qISL5Teg/YIrMr7K3LL4uuxYwMJMsi5MmgzBfBFvf8LC7JItRtP78W/DZ
GCKD+NNlVUab2sJebZ1vnTatByGznsimYm0DU1THsKoI9HAPl+MQ2Ni4kzd737f31Lapzc26KB5/
imGHn3G+gHT6y77ZUGjsOLwW5U3kGmQgUsW62I1r/+KqbR1an3nkFSMVKKVIaIVBiZBDt9WX/yBE
cqUnR539EwrbbmDz+FQr8wI6/RsT/++P9FvNo/5UwEdUNCMdBZgROjv1M9K0ML2yZtMlpDxkmz4B
F2+Svx1+VX5u8CBJ574+Ue929tdamu7aZv6UDF8i7GigHUo+hoZkDfPNdZOlPlLYLNZBLszuWezf
QaHzaLFo9bKoCJX++Y5pCR1OFPXCqK8EsP6RqmT0L8AlCNNtdo4AYv2FV8LgddOASu6pGepo0E4O
sT965nxWjsabze7OorsPIVHJM7H5GyOXmjTumyqNGNkG5y1zYi29PM/w5wRrnOx/yVDHSXBxFG7R
a6TxXRm9g4sVc2ZssLPNG2TD+BgumU2dB4YSTnbk97GRXUsFKFTrjVQ8fx/wSxjbtbvvZBvw4gjX
K5tI2QzjKQQkWJJZStKTG3gLY6DcHg+ho4ojN6mIILcp/AYViXaz1Q0WxJSp9/CfTYeHQYutw4Jn
q4FtzU3Di5c0Nzm1t4wPHZxr7AJCes+r2CqjWd7hlyeM4wP+pEfq5yTYsqIXi3mOkLu4swZxVHiz
fmUr8rrJbKI35P7UYC//mO7QtUEpkEnjgDO+yk00vUlQAI8tM7CceEYw236gQrq4A6DCKLyIyjBK
OEnd/ulkRnrd9ZF3K4wtZST1rdHuUh2XL1koQTH9qbNcreyEUmK9BECP6s+SeY6WABA5gEYsBPx6
SQwXzOzEQ/4se8mmxHdNUXXzwzDMPWQeIwSvy/UX+tq6qE871kaedBFL9VzSTmMLc6mtDyDOqMnP
rdNiZY+m5rYJiG/M/KOxpFQFG51QkW0kmWW81r28FlhaRG3wnWdV3HRLj34Fbs5FcpAPbdLlodRF
wP9hjpXe8KCEDKnuTHWHc/sEhND7lWPCsJjYWNbuveko+5zEHpsEbH6B2YEdLTPnji2xFgpkGKkO
lvgT9EJ4FHEFsbQheEAwhWtVp7UOblxJBVm6gXim15/iSA3qAasGn+DNprl28YgFOlNuBlOfe+hr
NtwDmMbECs+Aj7fVcAqcvitVnOMFabbzrIHw+gm/5hhMMX5UhOHQ4y1FikGZvh2ajLXmvQ9q2WtI
Q6TdB8bwt6YqBoEvBqgFBvg2EasCi8q4SCiDcUFnblsH14CoH9ssI2vKqEDKW7fxwamboZGF83AW
qFZ8+KL1hEpg+byG2MZINMurenwUDlFJQ8oxDhJLbhb1FpuO0vkC8tE86rUGa7TFPfa/RB4t7b3X
ZuLgagGMjnoN4UJ2eqMLyK4Y3wBNru9D5n26qaayIlf9SMgJY4cYwbyG/p9ztqhmiEGFqmEV90SS
Izn8V9vSCClXCgkljRgoUTNNJRmgvNIzZiIluwdxOn5JZu6H/n3+wTDgZe6qp1hrFmOGDEmorZXC
EF1cDSGUCYAAYBXOpZkfXyI7nl98CtfLHXfBcf56GPiMb4kHdOj57tWSJsODcQrp55HOJsuVaTVl
oRMcY18qPfMCFbLOzCXPWUawb5rImxT4NH8CsE+eJTq8kg6ZRBr4TrYxJWhMY5JwjTCHEEC1ZN4C
4HoTAHClMKrSN38JNAXAJKlFHZHtrQ9HhXAeeyV/GC+6DZcp5I2yR4Fl7wz8HmHpdAaS+4wtzO3F
YudWgGlkpkWNoRieZ6uvrXVke2/ZPzMt8AiaGAIb4XEAcaSKUyi5AOiXxTO8qE5Lyp7rh4kdApS8
0HPzlBRTqomTbFGW8ORcwQ2pPXCNRPuVXyYiRcJRmx1TpCGXve5bONd1ppcQwfvJNA5+2vJRzbtE
t6RtnVziV8ih5rkbmTK7u7OcM4lt8yiiQBxxvWmIBEHSKug69qZB8HqvbH6ibf8JdFVZG+iijqcc
TX/ZaJpEfnJ1G8Az/elHEv1UhAjx0mA66vqyCcQS6rezHlk5dncj7r89Agom4S7zX305PwaxWJod
Hmv+nAcQ11aSL65KcGaERoyz7w6nCEvCk71YbqtMcmipvV2CSgKSTGHugQBd+AG0BFALoj0v446j
MHqQ97DvznazRPaqjr9XFwVlZOoaZDCg+1r5RANFxs7VgI50oXKmdhlY3CKbtdb5t12LGT/4OlOW
Qlfv/f7jV81rrbEbriR1R4FIsYBEavt/PxzBYtpBxuBY+QL7/LrrthhyRJ87pnVH8rlP+xvPojIE
4Jdn2A+Haug4TweyH+O9ZZYiPUBTH+fGlFq/Qyl39G0AfZyN4iiYNxoNLKDqhzBsfRZX3gEAWumk
jm5+v/+2lOrgcqGSTDMb9LfYIaXOXD900NwZ4tY6Z7hRys9kSr3HnnXtP+CB+p9rdmntCAwNWZc8
YHOQYvsqXNy/TrmygKizREaitGfebnk3V+LrB/YKalnYDX6nfJv8hnyeORS9UxaCcbd+rWS3THmE
S4sfSIZSBHX0lhMJASnh0dbzwJMlRL2jb/8liUxPZtSICd0HP6M6trQjZ1Svhol5n+IK2cxWlnDW
NZoyjdLb8pivHAGX9+epAUDkY7Q0UIFRZ4o4dXrvB/dJht8mrHDWOOHhTJrbkz4I2YyYINYjxIx9
0+a8e/tfkBISla9DCT8jTM1kg73SW6WGv2NOq+Ja3WvTD3KY6ugQ0ApWHsA+RWnWZn7qw75y3XCs
ybeCrFzTROgF9rugmUWisHTIAjLf1Crht1/cNK4JLyZ8BYwuETOSoIzRC14awtwvAVhItYT/pB6Z
qiQAqfv1RqQvTufto9AQevPgrw+mDFJjLCwS+4rVuRHhz1chz0HKMEqLm1XquxNnus37jcZyoLT1
ZXIn6IfG1WncvYKY3+0aCRlCzAmfODMv5c07H+RUUxKWc+143yMqbvQt4PAA/7fMg6iZzefKJyAs
aoqD+ASHavBcmkgaaEgyYsaIgyhCMJzPdYGFctazCV5VGMkvrrPbkn2HhebGz8KNyOsEDhFcF2dH
v7wzHwuf9vODDHTorWIBNlQF0lv/ruRP60lF24MhkfkDe2ZDDJhl2O2OOQGeV2CKu6AVsh5rJMg+
earYQ9+O0gLGf2P+BPhTDhEUVc5q6mzPSnqwsjhnqgOg0VQSuLEC6rFuYkNx0jeQUof0vcTpC/qU
O/EfzLpg0I0Z8tvYvB2TYeBB1fbZZ6EcP0/XA7btY7VKkH/nmtH3JNYBxsAhsXCJZ69XGYFIME0F
R368PGbBO5KDE7GQVHe1dw71Zz7AcBUQ41jGGXmHmj1kHsBX+limEdTgr3XHzQRyKJhpcC7WJTcI
LZDq1mNOSbsDXJFYU92XApKtNAYjC7Dn4LsHpGjE89R6cBvDSWKFhU7MBIQPb6mcp8Z+JYpYzRsx
wLBqxzjvTY6jFaLJ3EQLO6ZqfxrbxjVopRxKFfqKpo3vdX9G5Zvx6BeyhRpJaFva1ma9vsJVFEI3
ZK+/zqKBmPx9A0gbJ6TmVlqePk2+JXWnSLas+5hiRXVsZYtusGQTWvBUN1j6RaPu3tkRXqddiyah
LjPTaQBNIXtFqbOUBYLWf5A4InKwvYdhP+Ewhii6dE+aFOX83MA7hVpbcCIJ+ps2ehruK7ZAs5G4
7KZC2Its4mdlnQPT8p3udXAOd0bd3yQw+6pekh/cXMnYmnGzLfKaNKZUDm8xtxmu7e8jNGXF0cIg
iVFBHPovc1oeV1BN+nPQMoPMxOo+jynPVqS/MpS6oMfyilUpEd8QFA1vPGRB9s5xo3tUi0xdgFpf
gjWrY4kDJCwVB0gpiiml023kFr2qd0oEuNtHzw9NYvnrhutyf3LsUED2qVgyI0ZmlfQHPLntRO76
TUExqatuABM1hifuh/qM8HUnn+Id1T/vcHO7JD4w37FSzCkx78LsMnevegCO1foyDoNo1Pi/aGgl
hpy6Pn1VtTA+3bK8mZXo89clRkFOAWv7/ZHM3B+UL4x0gxJmRfnGxXlFjj56hFM8eIAU/PRkeuzo
XBpFNV/EK/277c5WibBL2vmTWKT3QttyGWPmed8OxoSR3b8k5lW3FeOmfYvFyR1cFMHdRptlvOOx
iwjs+y2gMxjckaXRenM41+cExdBMHa+ddCX4MNDLnV/55KpLt9USJyS4a39QZnvS1lqErGnPOtfk
0i0MHmabSUkRdQBie/lmwhGIRqTBKeoMAQ5jESasSEYG87c++DYH4HNhRZSd5H2ArPsTuqKt/ZAT
wSPwNtvh5+kqwHPfd6sART1ZmwqXRVOtF6y2jRAWAEvFKDar8PbNvxuY/irBuRtdwEJYD03rBXvu
87kIUBaoJCz7ksfvEy+rBU2gdLyZq+ihsACSsRKD9rtFn878H8Ysf0ywvjENmVBO33Oog7HGf5OR
v5nLJTnlteqmWhxvXt2O617bAjPMYzkbqocKwkqC70w0rX/tE7mR8O/SH7DIYzGWBV/XMelJv2RQ
nkL8TRSiDfqHG2L1oxHcedI/ysvQW9SFomKV3ES1uiWDpjpBGswfQhgXugkBUNGOFrbFPQG3P151
esGdi2ayg5HZZwTTOYn9RjkawsONrAl8mFJ4FQDfHdqmlbWeGd6UlpHqnnNj7u5jdIzH+CbmQsm8
uKBX+SF8XetddDM5sGd1K5Odwut84XUaLv8mmFvJPI/qrTOCgnRS6yd5QGrR0ztsuUj8rPqoIxJW
yb1ZENobcnGrmVlCLeN48hnVCO9Izzk0fP7tuddsFuoBsXBM5HroKziX2qRTZ7dfLIjfXPn+NcAr
fZRvM6R8+pZkJfyDcgk6BCQIOh5hlQSSHM3nsGNlh9lHBqVWPocHD8fzOmOyF9qhG43/ruLoNfiL
3kGc1PuFCV3w0QT5fGUTVXf0LSOoyDS/oP51gOP+x+5lfE1Fs+IVF+3Z/0rv28rFFsdus1i31Q7h
CDWDWaYP/PbM3BT5Sgy7NuO0CI/Qh08dxDb0qZI3VAiE9GNj7xHGvsAiFGa+yN2VkdvvbuGZ2cYU
jJuN4WRbH4gwyQRY9CV7O04N7c89OnRNjValPQvyuXCWWm7RGYok2XeY9jnWQEjR4VXbM9G0sFgn
2OKRe6yK7kd3A/tU5qgYf2lLUlN49Te7kl3CViqoQyQR2+2bHTncK/O5mRM+GKP3KYsgCrVYvrng
MJZwO9iL6c+H4OCIndV6GpYqJFEqh+zcVeci8WkyRZYXdCPXHq9J1Pn8jYXVK022WspiFvt6pesd
UnfM+t3MzTRrtTdwIw55Dqne+Wp01COZEKiWtWIsC0+R+Mk2hWwswCXC7Ld+LmV8w3zLNsiVcIqB
LEhD4VO/M+VKNgtLTGM1mcDJxMetosrgR6lgYlaY4zCxLOp2gCR91q6RnZNCeV0zIbOgsvH/qqQt
l8dlGqpfJ5WejdH8Q3nke8F+vz4+P498IGQs3q4aqVf8q0tpYAOXIHXyyB3Gk46OMCfXPTY46T/I
CinR06VW6QT0OD+BX3X/r8zuMh4cTbShBPY9yrX3m7Lig5r6rCR4x4YtfkPwBI7xbMmZQpxIYAfW
tklSpPTxrXW4Tx2l1ShsLcRwtrQ0lVnprLwGt/70YXcv1Ac+FvT1ESl9Gg7S49MwdUm4a5/+8P/l
sqOBKp2gFnDz64QTzIguzh3kPlvET+J8yGGczpJB9FpEm9nmC7+VOEWnnHWfqqBzi9IT4UEnu4RR
ItndIrMQGqCgAbgcebntga/AFM7t312rVCkcWu0gr2ZGXOE/67inQHPh2LVtcDmN6Gl3rIHUkv2x
yG8+nwS+gL26jgen+BB6Zk2uvxL8BMTV8wa3SGSVweYGvUfUnQCvgoLhZHezHToREjIh8n8TO2dy
dnkLszP6pZWTlKCAGjMaapPZttEOrG8ee5SVBhfOGdKrzNAcODcsl7FCO3/amAzjL0uYKtmiIY7s
p4voKXutnLJ235B8PMbaM9EMQSdc/eOEYFZR1B4g6pMt1NScJtIX0Di+w0AY+t1ePPRa7ovJXY6n
eQbcrNFGORSVvAFGI/KopQZNpxQalFjRAOplnA2mpdIukajvsAcTf8+T8WQTdnSTt8STSw62cf9c
BaQqx++IvdFlGevyDkx7X9sbMdrvNqoOhCpqnCvyj8As5Y56X+agsOUv40tsHFK74vQxnAzcUwAo
kZRXl1ozBrCUKOkNF1vf0FHnZLwFUNkDd1e4BLEvnaKQCow5BEww+TKUsZpcoW9SQyvrJCqLTDdW
d8lKlXJtUUNPHJSABaJEaM3QOnm4SY3JEBPIZUY83+pTZ8uxgeFs5Ob+r9nMJWglrhQ2YoWcHCRc
XA6JEBoN6KdCc1glacB86pd2m23qg4CeIyviHDcuCaKBReEZ8hVaYyZMMovcsC7x7grqPCJmWv/K
Qho6Ly4tO/53/pLGXcpsgCLID1WtGI38LbXNFZ0didxJiv9i3PzXL9IeXmECDfa3oFEvwdl+CU2X
Acd7ahLJWsE0CM5iT9i4hOvD0C3ZdcqSmdfLZIYSDqujwSu5c3z/3Kr3kkU/RYQC8CcaB7mKt7JJ
k8XSZpQ3/RSBng/mwZs9QFkUUxmwwHaFSzfBXxNm1t2qYAsTPCu1yDq3dURb5jWnYW75K3/EksbM
2Iel6Tp8fff8HVaeS+n4cCZIbAjhNoE0ZRk+X/l2oyPsHeucWo0cf7vUYxAFg3hRrExJ8CsyRgtR
7V7CB0hrSQeTEXkuS/2Lq6ryMgwRPGXjhe5Cmq3w60PdOLRzc6gpKLNWRoxjp1wu8J02KEn8ajWd
Rlh3BEz+W9ifYb//4pt9lhfAzZyofVpNjijxJKkOjUQdKWg+t57xs+ctsyqTAiMxPzsXqpmMmnVz
d2v1ypoAuk+M6gCWkuK8vP8bbXDJLOfkJJAKhUMp52nxeL7coT4eUoACgf9Uv3eVSGz8Tl2KCJgU
Vt//a7VnmRJF9V096IWxk+YnzQoZvIhrfgi1DUf8TBCvpHHP3CNK0XnbU8pmKguTijPo8JaRAY5G
qrLBYWrTtabeL+GakRcPBpuzBtu+eqZRQREMpWbY+wSMis6EFQFHee62Hpa12KFOXQLn3AAgXSAr
+4eeSK3Qt8iob6f7GPDdDWQ2cQjM1237bEIxQmtxDhLaKf1X9Jp74/7PEOD7/a9ZuM3zmV8axOG0
QQQ/VnleEih8LbtW1J3jKezAor0Yw4mD31EfowBLLcD9vrXC5M4VNiNIMvpQYzGtHkN89rIOz4cz
7DnrngvNAPQ+5yoO5SYiOz/Q6YJgeljkmU1qteZJRJeId5K/PEQjDfUEfVEF6ig/gpSPyfzNtKQd
Y8ZdbDEM21PpwD/EtXzIRsCfdrFrjAd5llvqQXEGvVfaf+Sqw8rYwRoCeVzuSGyXUx6EiFi2tbC4
0Ka+O2TX8R191sfrMhTApMsdRmTAUcip3aEfZhSnVuTgUd2PfXa5hQJhClcM7Kub1e3177zlaOyk
am/D3fWo+0NktlGijDBFh/UmtnBohDyrK4DzmzPm5LmknVEDV2zfVjN6EP9U6Soa808Ym0gnVWqH
bA8UMsHsf6PNQPebh2BNyd0jEcjCDR6JkD5yFrL500q8hqcw/La7wgmhSHEiuHBYObC7gRX0vGJ0
WyaREtfgs+GKHhooVyCEinfDTinURW4rZnTsfCQmNSYPxI5ELQfdfUlMdyn21UlFTu5BmJ5IQQZi
2xWUrQASnRPffS3YCPp0efoDbwYP8bYmzqn6nTd2r/LsoCPaO5Eg3IiD7XyXnWPxsThv0sUJInYJ
BJnUzptLs0zsIBXV+J6EvA3CaCwZ0Pk1xPh5J6Gvcyap2YLr/SEJVQLnw7RRWsk7uKlShocPNBNQ
m1m/uIORJUMicPSjyHyzcb2qyKe5XJbsTUKOMlCC737GQgjB1EjySXcYy+XTlmk2tqHAIrJ7pTo1
1egTl0lHQmOSXru//ZODZwAdL1x/27yeTpZ98viU3dpvwEpvXP6dp3nh5C08j1HCvJAthfE2cSK9
2CsiqRfHNfVCEdlneHaUpKY9K+wNaU7tKTiNZfrAA/nwVyTLmlKtJ/7mB6eIaYs6bvPgvIOxZGa0
XySvS6pUIsS/cYdEXpT343EqVayi10/1VkJjLzWkPg6kRjEpPz2+eC/gD6k7uV0ms9Xk3tvQaIHF
l7lMiPDTXy2XOwjRQJSFHFF1sJ+qtA+M7byo+djo2zyMltlCG5sad6nh2+Vsi9haSwwQLGF2esYx
sOpmajTE0dbGIzNoon49UwFngkEJepcdi6laicsvS0dy65qauUlVWYSVVFE5aBb2GnI1G1iEfDlo
mlkyjeS+N0ZNRglRXzSBHwLDt1KDDMgepJyteTzJ86rtG/YjIFgYEoLE00OHxs3tXMDFX++TSn81
x8MP+9cs5DxLi9WH2khgoIuiOoCX0G730ArzG+/T69rBmp5VxEaOfUc8hqZZAUv4DQCcJdwRu2Mn
2r6ej6Fv9+sWxsnY0BSWyH7MMiUxnzkXDo2rUgrXOaaqPGGY9F4Qr8rnN5HDdE8LuTeKa+V4Lack
FmU6OL4ZvN6V7f4M8XsNOizcuu5BKWcFO3peKXOamtJNccDoqY1u1k4nWk1FNZ2TeliwpXZjuvB2
fXJ2ULiIdwjCY+Nyp+fXFJnxeQOR6QWkKONmygOAN7WBl7uO17vF8vKUzCAe0Psz0d0u1WP4GCt3
KbWO3gNvaZd7UPx0u1kgrnoBr6NDsxzc0k58g6Jau2vnkpcajX6oyWAJZJ6I5263jlt0N8eB8KgR
KdS9d9Qd1nf1hDI/biwPwCOgxNn85BPCDOFKh1hdwT3Lmze/YVAxtrfEMpgVD7mqF+aYldvW0E9k
mohjcwnKdVs8/2IIy0i8pLtmXWhI/LiBsv7lSDN5VhnjxFDoe2RBGhFCpLTMKgpPBMQCYOKQD4u4
PG8CnhiDSTkWjqleW8LyqpyoRRQQbyPU99SmKPwuUey13O05Os86wkBlL++9RbFLXezF0xk4DcUp
upidNkwnP3LtZYuG22iYUikefuvpSi1x5r4+ZdhY6lWlgKGjLLt2JYHQFYjxTBLaQ7f2UoxQYzQD
reBhaQcdu8xZahek/RHVP2/2hCeuwxC67bcrv1JYSNRalHet0NhcVWfUXmVcECNnVBZN2cubkLVX
o9PGZbmIXY+YgR/Te3ET7H7BBPThRwFlLgDOIPDhz0mDzPphg1CiTjWyobF8eB7XsMQ5eu1HTfl4
yntigoO2+o/W60v/sHUmC3B6rOLrhJWazj4M1iEYIg3720KXCJTheohxL/gk1FZuhzmbR8dIaxy6
0HUKGJ0EBVr9x2BktdgNKlQ1krEdNhwbiUYLCyaoEv19Qmdw3/I1mLF3yc95pgSCJqVMrKHuwJMG
QiKkL5JSXQwksZZoLhlbfkj0amE0FJf4sOhdOIoKka6MOU4m45FHHIE9DqzTaA20Igor1kg5x/VF
dx6yBdw1NS5s1SU3/CTqNbErF+k6XpDcAywAi3ud3tXDgGkttF+AcBXthyLFr9QuKRXjcaAamkwO
DLDYu2kmS3BYlmTQSFe2z+Bo1+LmBbrnFKpEZPD3D9qZPrHS262XL5dVA1LP78ILEkJ715Ir9zuO
bcjUsjb4zsUPu3zyojkLZiZtypkUMqmyvQ2W3Q/CLXh3Nj7J7pxU/hSY0+TXhxIVU5ktSJ9M9m52
mRPVJvjYTh1XhZygy7HNgDe4+y/iYMhdUFEM4LpG7RTdAR+TEYk62zARXtDxuDVh+O3OiRshQPlL
UXLv61TXPtGrwMwWpmHfLT2bMTH2quNxzPjzY/OiAvLjhxb7W4+IJeF8UhP8k+4ULIWtgnve94jm
A+koaenw300JbiVblofmhbJ0LWoutpfgkGLS1X+C0t9rl8Vm0gJ3lxbMP98o9/nEmeRBGIOweYtf
aovMTWQa9b6sQPp5iU2iRufL0WZnbhS6FifCwaNxDbDftVuQFOoiPDVLAb/y8KmnNeAcZuVVDEqY
swdbEZNXkDnaOZRiU36QbmVTa1BuJ/az8PT3fkF9CKyWjGUYuDiycbaZliPRtpV06OV84IxB7yjB
5qPllSm9aQPdo4QN3ns9T3Rqrr81hek/CYNzbmV8ImWvtf1gdumiJ5IsHDV6ZDuvM8xvQWTJIWWW
VICY2xdgVJldck27k7PZ00BQhiB/CWo1W9A9Zi9iz1o34TXl3HbNB15vmD3BzufWsiJsYJuW9t0d
lXhdnZB9u9PWypmCGf//2Vu2IBYFUQLL24688/JQCZ6B9/qSViBR3Ad4tGxYVEx8beNIIwCiSuHf
+oQlN3BSrObCWOV94eCYM0r8pw4ROyCPd95ggRJjVarV2DjK8QMhNXq5j/97Q5J9VMkFS/jiFDBk
0pIZTXWdS+/fblHuX61y5W4VZTGO0GNxfl+eAzQqh4J/3ZOTSn6JVj1aNZbP/IIibdyHriy9lQLD
+aWxbjUfgjd3v4vVJ0B2fHCgccfMayHAYXvrwiMfAE9aSW4hhRH8aqDrO8uRuo+Z4BOxPYUC+0yY
e0GUZSenrgnSQboGrL8wd3Pj1/k8u1QBWcaVfIuO/93VYUDr4EXLXe+bfxvhdLLNS8bNWNoEvZg1
s998hlc1xNaXbMWUOJNsgJz7tXr9/kpR2L1OjjX+Re5+tKtGiNyH5KNP5sDFzdU+lk2AEczQzJ1b
RnEX+gDQXSpca0bvWfpsuU16R1AQ5WYvl7urULotkBtuJhJpK/KmJrfctu6ZPTJCSD7HuXNbTUCh
syPSd3NFvnDrY+/7bXRF48EW5OfojzhGR/o5AaeRqQq6AYfiLPCK+8mKrhFyAKoVHX1vhEEgwZ9y
osjmhq3RKV8S+1OogPEyJTp5ODvrnBMXYvVA8Z130eTEontc2NSwUCp2xZpRMVZHEpmXLmvQTU+M
Nwv7yFspgih6H0xpo6wtal9MW8C1wdpqJkbUf3jfQIB23gAc9qi2RaBqZKn1nyYcNe/QFtOr5w+G
J2ASCtTx59cDdQ+djoaKHuSEJVgwXc2VHKX8h/XrdXsOF/gEC1uPP+6ok7sNaBpGvdXPjolHq4SR
0cA3i473O2rd2iZm7oceSs/0at/soVbh7NyVjOR983dIHh3MG3O/LttrPaMugPXiB7bNnWFIeDWL
+G47H41hZnX/oVeFYiIO4B+X72Vn4GdQ+B7uXGFH/iP5VoDPoZjBzlSrhcSH2eqiAwd1dxVS5ans
chUC1LUO+VByV5gnYOovnv3jQPXc3qs5q2vMtWdlQrebrIIN83c6OfdCo+sXGhLCXht+xKnUByH7
ZaF58VApJmIiaLW5a6C7II38jwIOFczjPcUhM0yvuzxELTES7077MPuEfG1mQ7f+XajXKbjErHc2
KA9cSNtT9zYnyhL3IJua3e70cSuAF32VmQvDaJRQFv92sZxS/wfu4IHiGtndLIVaDhvFg2fXUi1d
DGL/akCjOPdCB/4Pxf2/vCxzqhwen81lB/sHaTBVZl48kna83u28ALxnQEapxNMwwzkqWr6PZwVJ
jnXbr1jhPopTJFk+NlA8Mzt9X1ahkrDPfu8oYpOonjvvVMVWXA7i3dI78Prte9C/UyiYHWHjBGWI
cferSGnVl3wub5WB0OKmxifMw2r4GMNumprh7+CiiJHxVwkcgGUKtF8MtErOghSHqQf5gKuGwpma
OOzLOibZh1i5F2gPuHmKV7Hk9tAoos/df2FqAdV4AMBb9w3HJkQ0M4SI1/kbrs2+PcEsWZMfgvrs
svY5xBoONlFAYS8a+3OvZILepzTqdPuLMBUdN2XJI+gPm9ihKns2fPgjqs4cI/H0hVzB4WXwqkEn
62Twvd31MUQNqt9n7KCosAD3jyykPzvHNLg5twad1YXaRraXaDSp9RZAb7AbInwDs/iA32f1JvDF
mIcotTuQldJv7UAb91sIsgXE2jhCIKZAV5gq91xSCvqvSMGTN2/nBUmHb6afQM85rb1JhWj9umjJ
sCkzSqrr73GB4bHUwgNngeOWzLgUueZMmdk4DJ5vvAWoqAwIE9VG5cnnfGkgUF8P7eq8ue9+p48b
2TCx9wHHFTbMYsAFkGxeXdnph4FBqARUqokWaxw/JX+F7IFehNYw9iRP5qw+nCU1Q1TgeYPzztzn
5CTeRjieK0RFGNqXKkvkxA5l7leZU4E8wvACoVAZlDpTk5oEa7nDj7pYyVMSp8Q6aInLiU3CF3W/
h1WH+3HvizTwaKSl3WUNJWaMX+NosSzZ+8E2M1bFnSesqMbO6X6UGal9xW0KSUgUbdumj6CUJR6g
km9qmuNV+4zPO7eeFgvUwNkCB1DAfYjSHtRCwvE6Rg/IrsKry4oZ46cVt48y3f9ApW8Y5ySjoHI6
tys81G0vjKHk3sh//4DOJWoGFkwHE0kYkK4u+exfKpTdSKXn0OE1C0UcSYVEb0rgEM10lPNjxd/v
Zw1isbiHrlPogY7R5J+7R0ejGE+pwKtnou33yuVY1QlHeo2zg2AhBC2LPPWsEzBq8OBrDXgbsnIJ
9Mp/XZGNLBHtQPZ+c8ekmBbQvTKMsbbfI0oAdUm/tpXPXHojYkHrR2qxQjnrwLW23d56vZQNF3M0
lrO02JOsQBf1y8/Ud3v1IiYKn3H/IYlissDbPmv/vBuYSYjdBftZJSX7msxJZN+jiFxEG2j+RX+a
U/SbbFXE69awl/S3jD2hh7nLnt53TAQnJxMk7fG3GYCUiEFCGo7feGV6TSrZM6L+brkjHnz3eF6M
qvqAY5UYG9oz2SIRK2j9lz2uMP79EJZHeFp/mwQYCYy85UXVg88io/r1Mvzheb1RweDOLU+FILVH
fBaJYdKl0KOVBPwcmfk0vbldDtWXgP6XQZoM5n7AxYMrsirdpLGIRsjnQqZbWeTnWLz4D1AmEKEn
LQMZHNKqK4NwVpPUQiAyr5HO0zklzjv49UW9bwyR6SpT1F2N1w14Ldd9VMiARNhqAfyI3Q14AbvD
VWXlmPoEaVpnf6FDd6dr1DnXra55Acz4QKpMdcx4UymT7lolx7f3lGGbSl7ssCTB/ySzkVBcuZPs
uNA9yG+ytbMdZ5Gg/TA7+PKNOJ8ggf5ULTh7OpYOEuY+o1/mvFWBLO1nAV9YPq+nruyVDQpJW2rc
q0JuM+NHqTBpAbcZVPxSE3a2b7ZsAtVOhlrrzGomb0nTVmROwytZmeEWqLX//+8RdCS3XQflIyKj
YFuVR7ySyLu3FhnRHqXFm19Bx/rvQW1asVwqeg25OPn+n2AI6oqS9Sw2OCTwEJMzo13ZLoOo8+ua
lr8Cn3j2ZGxzlzySsa5rb4lIS7KXCrKJgu6PPz9Yo6rx7OKY4aYzKa7ot3STLPpzP+HjsmlmpL6r
bk7mnqSDmBGONnWODvZej3HzM3ggVDrxJJmpwR1qTdWvZAVbqTviaGFowE0mNqpye1CGbGPlquDs
oWeVvRxZzApIcfnYmt38X5MwMc/M/pJD1X5jPZblsnPCx35am9ESn791eu0Mhd6UsPEvNSZ53tZv
KJG+MtGq+cHldcppqsAjP2OoE4cBTHJ2amIleh6/D1aV/Hm7Y9dHTkj70w/2vg4nB5vpIYKoPmuo
hOiZWMvZR5tVnNZZV0m7XzSctb5vYrFVylhMF/9tVpbDb6/7Y34RKCXj/i4g039eB4ZZgOKBePX6
Yr5YXr6RzrUmnNc5yV1ikmj9T6ZqyLrF3uTx3nt+lsnal1CzQ9PXV9g2ezt+55m2t6krQP4WJrQu
+WBSvfkhNt8bDxOzGaEB8QoF7BApInYaUMN7WupK88bSK2w7DhIZAyKS5s9ZbAwgD0kCzaybeLpm
8VFLsgZOZqIWggBk3/OLmFdUDTp1OzxuZOShBTkRgIf2kkJCOP2QlYYYErT9Eap8+oxVzuG8UAQ3
bmTWjY8oaeBa9u2TpsrExvnaHX8fqRHLmGaxxgYsgzn8Zqi5LOrpr+HxDM+wpRJ9/ELslKE68YPc
/LdYfir9jMtXXx1TBxBiN0VgOFDZHqTWJm8Hk0gKC9X6xC5Jb/OOyKjsDc7rckWhNKFOjNBnW2fE
4PgYRVgFAOLKleduZjUVsUCsZ3xlxRis1YEOYDXQ4gcdHo/bVlHTWLHTez0NrbSEPaz0klkz3kdi
fwHcA0V3YE8xKzuZUaP4o1WLiSmcRPGw9Qto0ij344olIh9I7pScX7qQXnXRXTgttFsxGLg5Mb48
50ksxdBW68w7e0+JZ/oqCqXXhK10mR+jSbqIWsZ88IKCaso2HOoBm/+UcFluthNCSVTwnMjDhK/5
pAJaTRdgcM6T0ANXAP0Q7Xd2Dx3MaxUibPC+t4a3gmihm3tNJMbk2ESbG9R/724A/CGUXA6ukS4D
XB1yMKQJAJc+olsRIH5l7ToO3p6hvYrPFMMt4wX/b/ZGBhhBlnM+R+Kja5LZ8QSm/AINrqCea+Ja
22RGNybx5yLrk5+ulhdMnc5iigAbG77WYc2GeVvTFrXMoeDRN7VIlB+7VyWZn55zxKdSuhTvNl3P
DZCShMZdWCJ8Il+6qegOqpVFHNinczIbanNv7oRSRItwtmDSDg8EtVSGorTa53Il7qHft3+9MStd
9jlsnNy5wR1ghRMM6SbX8d0aKs1AvnBR6JomQ8w9GJh4hP4YpuwL1IhwS9WRichsgodlJ8lNdZgW
yeMQiGaJUsMibN3kEyVdNTXK4BzY/Qsw/10pDo1FVglgP32kD08+a+VcAuL1ZXbG1pOX7/KVIMOT
rkBFOUXj+e0Q+Uyhy89iDMTIzKnYARv8Ri3kWpNC77/nFrQKA6HRefPNNMYY9G2a5l7ZszKT/Mbj
A5SHgrnS9OH13S0xgvRW1l7o9jk0LWXZs5UYjgGlPl8nWkJguP9UVgMEdQCHK7Rnd/D2b4c/npz8
eIX67nh+cpoTkcZGZnvHFvxF2itRmNfvjoLgKHpi0jUmArqpXdEttnRCxhEFOTaW0vXiBvn0yDWk
M/T5QKE7P1zx55Pam1cJTKgHibKprOoiIo1OO3TwxIyH7Ik7YkSY8CauF4bvGNAt4nGpZMmA3M2Y
9suGbqBlRMObdzRoUffDgqPNK+MB/KnHBDcMgw7liHiNlYnKDfUVydl5ZUD2KzWqM1bAGMDr6CT3
sK88fX/dDzre5CB+BCqsIzHfMRUvcfNYdZcjVYPlVaHum/GsYMo8bnaxC0rxCfpburRSEmrLWInc
e47xbQRbvzMHULdrKxFLovX4batpxKTIbQ+mpGA5WXj7RpkH5cKbE+bkgvY8faH/WdR8kgwW6oNT
6oPNqr2R0BFk4j4C50RpNNYnep58/FkONzI+8RiHwaCb+iF5faI6Fbf3rBHZGqcI+vQVbwweQweZ
RFHkqFpog1FxLf4TSpSzckqJuLT4KfKPItwb6vg7guo3cICuNIECo/iXDLyc52/FXC0PwWNQmmtg
Bc8TxW+BE0++nq8hxQX3NF2k2Sqc5TqszFbH4GAK8/1egV3OLsgopr7GYdWc7nlYEtTXuOQC1P7L
/tTexNTUw4jNxGr7SwNAqss88TOoyH3d59qUY11edJaRM+0Y8mL3dMYzBBRl38El+jJ8p9bLeCen
HFuwN7j7pu5YIDt6u2jj5nT4ij0caIBQ4nCP+3yxbFIBNV5dYt7Ub56M1qIVlv4lJzBmu+HXKW3e
t1haIMyDHGct+0zV4CVYhcqqaYEzkTN5hfbxVIezqAuTGe/ckVhGj7zMP55J/uj+00A4pnMvEHoR
kH6a5Lj6MDvNJXUI00wOyqLQCTRVMb6p3m4qDCDZELXsiXrwrEp9r+j0iubYmbaMLGYjZ0rwdYk1
Q+sC/y3S90NH9Qm914fGzF5ZUwsANoyuq+mW7aAgXMI6Uoz6m0Un0tT6LDWvhc6uDbOaNUmtRRut
QeastrwiQpnYAOoyezOz4dTAGh1K5COoGhlJ8Nx/TSe/cm3dwEIhLVTrl7UCVROPiXcyJ2krGa8G
TJXruF/BePWqgZVPALWAEVrcv3hWQG5yZolqCOjhuTBmjA0nKM/MKAa1FXSUplqh946Zkaa+1MlJ
Se2hIzaNkSqIf3P8yk4djfZCA2bx58eAJABxoOdpTtJYtCny4XDePDj67VmpycKvcRCI/3RKvx1x
scqNualmRzji8kOYfrIG16zBrfNr7cXIO0oBvUE2Km89hbRoScczuG3SOC8zRampxW+cCJ13STIl
YIUnLiObvHZDC4yM0psyXxcYy8zLmQ01ugw2oTmETqH7FGAKBmvSrLC4rWJSp29wlTthE9Vgt0Ox
h3xsg2hc1drGEDOqWPiBsiACbciXl1gwv0eZiqdP1mO8xjmA+wpdjK0G0C9leD9CFdv+50Ou9qNR
GImPVMnuzCiqPxBJ/mHZp2CVJMMuke6vAZLytnq9DSt1vk/U8tk37vCO85OJfRPL2d9Z+fjhpFMI
ZSqS0zKUq+nrg99ybCUmAfse4sBSDFUXRiof7laImFoDqjt0Nub07OLTJaKo7Ox5e3ezFPEzZc5u
mWNdxgNPvOMRLYONRbVKEbXVsusrEMJQgIGCiHwrg7YpnbvIqkbhQQhsJsHTubZdT4xwevucbpCA
Oj6pMIVQVP7zUiyiI/YylPgx/h1GXBY9oBoGZv9+UAo4iAFor3up1aa4NQr0SUe6SLdAED/P6TGL
lUFbNOv++xEIJEMBnbEYLdJgOsCzMWDQ/37+J5gg4eU/zHQn9WMhLkJ+F7JEMvIrv4gHRZSZT6+D
RQAfmDRbB1Jd5U1tcrI3AJj5Avd9IZAdgwezbdZl0FokzT+U1TlXOnFAHqb9Zy/+27BRuO8tamv7
eFLG45UtE46c8XkpSNvHVNtmiSU9iuXKMfnYqcWXf8EcdxSFt4xz4Klgk3YRV/o3J/tc3IYnjWwb
6J100pJdzmJdJuRNbrKHA7DS3D2thPnxXezH04kVlc7dySRBQW6xHCxLvF8UqGETOhL7B12W/Obd
TBwQQn+luZ/2ngjxkEH8lIIUf+dl9Ktl3CaSkqUQafwQ6y/87Pj/WocnuqL0XGmJo1D4D3ikMvON
2oiS5LvmZ5Ww5yu1lIStfjr0CVeGBKSwdHZUR3ziwk4CUa4G60yaJfCi/CJWcjzA64cCVAaZAapJ
3fC8gxShluwouvG01oggjQ6vSb1XwgUwJfZ/sdjk3WQUg2LKXOoHbNXSbLl/I/nNy62IzSBIspYp
mel9CiyYQXi1ZXoltbla/Twy9Kd84HpDMs/blsz8VyTkTNts0F9CrIUT8+4DR/7KD3mTo+3NBWfQ
5N0Vppr+hEbBy0AYeybqiBSmHWfrMG+fuUkc1hxJUUxe8L9o7YwpRVZFtARw7qz9aWryMJRcF1kO
++Mvryv/CltP7dB+7rWtYRPD5dd0toKGmWcNFBtC+EKEVYxkNtbe64of0jT5/2MLWaxQOygoSJ84
iJzbCeW70xPYsfxySrYKbJeSAwsVQm/VRfSENFy7FpPrNOI8pJO9nHPKnsomwrxrz2GNTHjdNDIJ
E2RzAR9BsI/o0PoWUApm+ROzMTrVVFv+1ElW0PnVUYI0V8ygqbK7WCPLfuE02+Plft8AB2vVs0RX
1eUiLgMTwHohLSKrZdZ/bA9W0tPF7nWHkJDTHcHIyDveeuhbenQJVv5B+8zR3+rcgMdttduM7yxG
CYM0fV6stcAz15ZyhShgdT++7Ew2RcG4R/bgODPdBFKwBB7XYS6OnxReEubGVjuZj3vZDm4ndzoj
d01ylP98Ha2u5yV7BpkkymmzGFt5E5FYgGAo7vnk6+BldBQyycB+MDcl4OWTPgeW8jiYcsdP7PJo
IMU5IfabIlogI+8+ptLQby+PIioVoq1Ofy/k+BrEBHOlIckDtOpc3X+UwYyUI0O+Iii6uD3iOPCe
Id29OmENvZpnJF7xH/5MMYqF90Dt4dEyjznKFd/AZdG+71dprHylarF9+/5Nj3WB+YjIlcay25tX
rkE6tnYgdaoaEqmcRHuew7bjHOqlyUoJ3rcg4mm9ut2MEGXtG/kt91IZjGu7eU1dB177SIs3eQKs
PVYMWD4FKwXRCttWVQJni1bfVBoM4H6p9tq3ubbU/ApsnmfA7sM8FmHxHnfP4X7k+HaYKenaqCsQ
2fKHcEx3wH5DU09H9zrqFb3HGt2kSWl62V5pdPAhwfAxQpXfHfnqpCfjBVQvKnCt4byWBS5cWrY7
rC1XHqiePtvv9/8fQSgwEIBMN5MbXn+ymBuMBkwk1ZMiAS32WPsbqOqlmn+gMSrYQUmTBoQUFVd5
VDmMoUEoADZY5GeyGsDCeTx8LnVia7whr41lMu9p5MW2qNsESod+xmn0L12v0BiVCgbdJmMx29pt
P4pE3t/Ss5DTVDjNjmaZYU1Nnn5GajsHIYeaQ3H0j21Y9IT23HMjYb6ddSpwNw16tHjOCSbET/Fh
DVxytSKleA8G32PdK1xD0TWqN3DRPPcTp4uxmAjNHFPvud16ifQgEUDNKNu+cFAcN6i/r7MW3KXP
KHs04wRmglwH93Eo0HeBVxGuObh1jBKdnv1nKTymkwtoktXOsgCsUnE8o2FNDlmYQvFA4TEjaGti
WTMH9ebuV8gx/KNTyBhog/HudEBq3h4CIkE1516Gcm/IGvLeHuSKIFsKrmYI7UWvcixHNXzVt60x
owBJlBjZYGkuqDR9OKuvEOg8oXHPvufK1cMEQjQCq7JBtg6vSMFQ3TV93b6k3CMuiZh2k7TaLSrn
waMQ6fMV2ML5bj5x4voqyQhY+QAhk29z+wC9q6EYRhqav9yo2YMKRoch3LyZIsoSjCk5D3E+otWZ
jga8419QYfvpXOEWIpCT/I0VRUjxfjdAQ+oQzn33eWUDc3e4EvvESJbX/zS8TmdVQGj7T4KedyoC
O+e2itui8x2XwOnYtVr/peDPqFy1QIUG2ghCNoNomeHkOjgxOYaxnqU/51nP/bqYcDmirbXaXipT
//wIr2k1Dhc1A2daNwy/w0Mbtw57PQtzSRC6xED+kj/lP9O679ayAxYLPuRmvUPBrxSxGz+XojI9
p+2oEVlQuatR5TCt+0j7icT7mIhGAXV9T0DsjHHvoRjsEZ8TPaMtwS6vjD09VZ/TuSK/8H7X4rdF
4kQDZCz6LADS5kNF+dQCAJnU4h+vl7Pw3P5oO3mLPgTqw58xZqoSp271Fg5abGx5yK7xUi/3mIS4
5R9xGNf8plQYVlTa6lLqGQlPRKoz84O46R10itzcR28ViDR26SKyV5g61sd6oPSfbB9o7wtdU8iM
V2ktF+YKW6mJIGlWyceCxEHHlu0Y4e/bLVhxPlj5/e+QV8ZLopiavbBGvyAuqiRg93+EgDkzN8Ww
DPlv/780XJFyJGN9yvQ7+YnClk9tbHKI7N3i/97rwHY9maUPTW1WuJYhN60p/i2JWO9jf/9w6H5A
GH2RvKLL6NwP5hFbWsbK83Ul0yJ/DJJNYV7raU4KxgIL1YaZFbzEBkZ1eg6mE3r+MmYWM1vTQLDl
+kQd7uxqGAYbNqtqNaU8Rb1OyxU+nMvxVWeaDgmN9alXCRGsty7xis63zXxpcCy7WJMjFNnsv616
aDVJcKZ+k08MExUdC6CpOGGjc5KUo8XjD+bToXmRK9VRUQjyoijtlmqK2vMeV6VNoWFp7lxoCkjq
a54L8XGlTLWa8a1ezvBI4iO9FLFHBYWvvcf6fQvJNo5miZFxphRZnnV97ryOWgwjZvKDGQIJlpBQ
oDb+O7fPsBGv+WvAawFJRsP2sCqtTzQBxlNu478sJDLwNqeKPM9nV909+rQPkmsV7EB15L0ZAaP+
3nCTdrCWzSkCc5IV3Ut9nGIufs16WDuuSVY8IKM/G6FzYZ+BEwmCU9Ib7BeHqYkD5G75aHi3s9LA
U+bxlfiWyV9qZuVm1wOVXNlWHg37Mq7QornXDTe7qwmf6INHfOUZzAHGlNcMEb4a9R51GkgJTw2X
LvrBtin8W454R62GTv/ewc4Ci5oLYuBReTp8uN5i8DzoAvwSfuwFLTFej/TNncbYUM+SMTaEGCht
KymW72YcedEZf1NRm++INu55386FiwbC8Nufij3n0sdm0iITNCMy2UKo3eqi8MnrVW1kwgfNBCoG
Tj06djBLV3O5WtHcX5axZwcu4FPqNpHFFsGgjNdGqYc/NZ8tg/TtJP346FDqE9IOln3YAoFOjP3U
KPoZPFRhD/1W6BQp6+Z5dY8G95ciouskfxICEZGNB2O+LXEFI3c5LzgV4ujun8rT47W0K0vreT7R
9TVNte7fgHQEd3PsNHX5kxyuSWvEnwOgktnJEw6dgVnNdRhpeEPo7lbY9gjx2AZ5fmUmd0fl5Bnp
VeKO3o8sICSCRfMWic+Lhu1vDLxRV0R3hUKp/wyyNpzYNElUjn3K4f6CkvT1tkGZPuXFdSNtSdgQ
r7au2Qyk9BDvOJicED7hRxZ93PQj/jUsdrmNZOJgQYI9dibRM4yVW+iw2l91nsvf5fZos0AD9+PF
lS+D45MpfJ46WY7qnpYhqCUdX+ImPWuf6H/4UHI2gyrhy7dCMeuKTN9OpdC/Tx5XXWgmSvdCMzXL
Y8kHkyBJx6O3jwEQvWaCRZHM4Ayp2QSxBGmCAIV7vaQfiNtSgrBqq+LTb6The+eq7a65MpUDWq0F
Bmq/SIVIL1/smE9JMHaFyhKHEnefp+nfjLUYbctvTbocai/xJY21u+RfaDdrVlF0dFK4QEJZ9HNe
7VqirSUCOPCGkHnZrcLgw5cVSw/olJZfkgorAXoDtmuIiYW3bsGtEsFiTqj6Jn2HGW1Atys8pNYR
CnrxmjTG+o00rGVU7wq60JznG/g0JCGTNYt8o4hnaPlqFyT5hYgpMVRb0FUVFKsERxrcVrMRdwLc
a6kOhN+XH0tij1YyoSXru094GmkqD6HFL7OZf2IhPN1yf/MqCzS4Ge9OGBzPFJmRLPrZWEA3Nyfs
E+or+MpiaMH2Y8hNKkKcQMCA9s8oPT+Z0Un4Il3I9Y/1+pnMWbduO/qYVG2xsOlxG2EnEoCoeYAb
xIygsjcga6EAnE5OZMIMnTdoDNIuzeqP893bgOK9hXtjFxFwpSumulHmUOpct5eBPB36PhP4aMNm
+F5YRIMa1T4mLxWkvE1JytULnnnO2itjk7PNHpfqonoDizANm7bBuWPVeCWJtY4dfJ6zpN5eTdNS
cAWXd5qlM08yXUghBbh4k6BvELxulaZvoA4o/PixWDprPWplnMT+/y3aSSQVMheljEbfipr0TSJJ
o6lBOxoxr+UyzXG2oS7tG1XR1qXmmHFr/EiPkIt986Ts+HFaeh28WYAWlOaoLZcHXG04rpRWfXFO
3wddF7ew7PWchfB1WSyz2CHliP+7T5q+wEduhuYq8tZt9XH3hhLsXer6uORv3BY+APU86kwDqF2T
sVRAOQcOlx0EAG+NCMsvAk6OuCRNndzsx4YFn6a8qWPSp+hmkz2tYsB+yqR6FolkE4F5dyLU91S3
nQ1AdRNMAYn4PKWhqr9hgNs6c70Dhfqk/jcXig40U3yYFPanMcDGWG5iI+y5O1fKv0g/WX9BHlDw
EZL6fcTpysf+k8aYhln/8xtgdW8sCQbIseRJ1ejfxzfcqQar7dMGJkOTCiUJftnqZ32hS8kd0hpF
TsFWaj84PRTfv4j8/9HIXaP7pcFMRQTRTFwISE0o8SEgrAdTXFF/sf2ZLF+1qNlIfd0vevO35z7T
S6KDV24t0kV5kSjJHaslB7UconGwlYZhkRUhFfHaU2hqkTVUZmFK8RMObvojWRz1YxkuY2e5Dx8I
5LhaTqx0S0e4BmnZD+jdwN37UruRYfEvMCP7nXMd9paLQePI7LQQfW4ng1Z7J1yoOV37M3X3TQwI
b3zXgRZ/arCSb7SL5+V+1M+wIKoe6mtkTXZ8A8H2zVSE6iugxI2957BrPFDi2i10CvmOQxVX5i1q
SkW/jlIJgB5Sq1HAK4FEdPxc//ak7UPdGQi8spMl7FGEQ8TxNEE2IaleLSDA+jVhMaBfsEskz9Pp
19dxalXdWVpxVPlcJuPBMfI+1VEv5U/dAHp1AFg5lwS9EVU/zXFSFhYcaiY4eLVO+xgYAv59d3Ec
n33XMtvW44gLiJJNI/qYytGz10TGLgb0Byv81e3I4msxK9DKxoeIPSejUwdAFkouaoY9Hh2UxOlz
rFbiYD0wTOOogZmKMYVJ9a5MD/5kuNaEodtYS1lnCZ+04CD8XntAUZxxy5fUb89CsNuGXYaUnfUH
t6M98axHfks24NxyYaBCwDILq71XJl780g2VbevDAItEsBWTULARMygoKSUMeqSaJm+V/cTjpyOj
uaKpMfq8VS1SV4sPqbRTL7W8i8xj1k6B7GVYWLm4r3djuicRHW1wmxeRlFVvggw7ViA1i6Gv0XOP
4xvF+QuPzPKyK+wNVWaYvCvbvmhT8GcZph0drAJEbMcLSiMdF9WayX53YNQjT3MJfFS48YbfaBaj
69wDvZ3FRLE9iYN38GvIO6qEK8Op/ZhHcTWirTjUaDatgWssBORTdFCEsvX0xEcxX+q06CSbu2HC
EiPeIXl98VZ2N4R34OgWl7wdvb4z5hCwecQzJUU6UU/JvaNilxG7fJ8hj40Lug0Gxx2BV5xVFZA/
i0Xxhv362NbsndWm9tqhvSv1PIekIBe/qmH3H3RRnThIOqWxcSpOBRnflvKyMoLtdw+4S3Z8CBcd
MxG8CxurJcQ42o3H8nT/ABf/hTEl1C81FmyjfBgWqAVYZS6cZIjLqDGyTKDohVJjUHzWG+w+8e0K
t/S+rGaSyqpBVLscEqhUfMVC7dxgZKgYI1qS6ZKbQFU67jJZHsgFHcFS5rsrkvneGug9e/hLbVo+
IrtYRlAYUC8qK993j1p1zKpb6r6e9a1e4/Ij5uzGXkCe0r/k4Flku5U0jeU+hNqau5seJ/V5cpfA
5Z+7p47zmAI/QY55BLP500pxEcOBAAn/VJqM/wqo9gYZTQNdZujprmQMgJtxQYT+nDP/t8wLQsOu
BBd4+g7FOB3oBMM0jET9pBH6At1vTeuOIPs8CDtyUlZQexTTmNm7ZTNMF4mhu1QOF1GWRRbYgWLE
qh+ynKP67y95upTwm7wk8mybLnJ5xDRZMBbtwIu9dmQsNuRhChhMHfP3pMs/MQi/wEZ+9q9P5iYa
jm5f1OqyqpIuzcDBbiJROH67UDUmA38ZB61l8IN7cnCJn3Bgw3eKwuONwLHBWJ9P7I/JBYCw4QBX
qbLsvJyqzpbPTCVmwCNNja9mrOhlx1meEiHxzgjW/muxA+1E3kwuodFD/yoHu9n5LEChW+H4Axel
jd+UmBF3xzUuXgO3A/wkYy6Oe6ypaLFtSJ0JVREyKCE3rWzk1UTc72LKWXQ7w8Un3WDC6rpW7zwv
A5riFcHHVgxmsDaOyqgPlS77m8vwKSQ5xSQASZTfba9C423tkzst2h8RtWA2dsUUh3PskAiUjBI2
wew9hiHIJFzguGK4Le8cxt1qwmCbPuBPSGkDDaN+/RaoFK5J/P8TgO2RI2pK9AOmeS2TsnMobkBn
HJZO9ZygjOwOaoxRz1U2CCaUa9baEjVvIHLFE/j1Y2uu5Z7BxCUsVOkEActJmu44sezO26bSV9w8
HCeC7Sgo1TRAu9LV3+QbfhEytPXbDUrkKhLU2uNJ0yDhQuRYVqjwv5qHQjvOyljF0iDc1v4Cze2Y
IyBkc4xS3xdewsxNXYLo5m8h517u+SiHD3NEB+52b4/dvhTyj09qgX+HWvRS6m9yn+dCpQba5R7i
1NEGXQb10i5DncQJEECQRcrQ24b3ItZqMeygwxKjvuEySVs6Gh9X+vJmeko4PiqcJNcw3lemmM8f
zZEcBckdvfZmaClbYPhVHQYzO2L91lCn7A7LRtb2QvYKVv7AGEWGynnJiiI8ykEDdNMgvqdGBe++
MOtyJZ1bblKan+UHXmo7n5xWqvSsCRDHC7oiYylc+Xy5ch41R5p0V9ovyqoZRTf1xpA1X5X667PF
toCbkuKUBILkmgNlAcxScaJhkffU5SOS4TyaqAukefGBXazymvxoyxxBMy2omDX0ujKgylF3fyjN
ZWVy0NqfCQ6D1R/ncsB+Vx+81spZqt0x0f+uDHk2WXjKEkkFclSpYhvO36SzibIpNYFNyr5tIEv8
vFGo8YNCjMyfIEGxyIPlTj8iadsMHzQVfzdNaT/tAV/khwe3QbEH5NJHXD9h8irFvzMdxd9rnnjE
N/7txTHkO0CaX7q8woqOnbQmpZLpbrlxLW3HcWVlkIz7eK3060ncKa/tPAA8yHM2QEuqA5dCsGbN
Hr17UoQyxz5AaNpf9zPvWpGRpmdRLzdNbIk/apw6cAIjIOKEVxViHTFvcnWP9A6d/yhWPtM3j0fb
XUkv9YhKfnvDL/Zvy6DOHMHUzTdulw/eE5LNUQ3AY6tZ9rA2WPKA1O2I4VlM/FazdXof+jvDxtR+
qYnSPMPszHkurLSKUt895M54uEounAmBMhxImW3dvfleiGxrpTr5r62v7nKq6/Q9txYXuvVJ/5UN
yyBHusAi01nWPHbEjar5t4OoKFz2WHz8BmraHzqUs9rXtkA3FOUIXkavs+Gmn+Ys4pDA1oEn+tZp
+b5Lu0bF5mUpk7BjP+3n7dl/VnV3aHs7U9yYxtTfdPiF7ce56BeZI+ulT7jqQi/TOL2JC/GkNIIx
pJrK8SLSRxopnjCxK1ssZ1hLKaSeCxmaiQvgIbza6rHBqPuEh1jpIPuF0EkA/DXfKqF5N+hm8NL+
uXDO5MYi+fVA6A5OPaddCV7b12UGuYOFvTSI8oDhOWLZ3NN4lpcaUUepignOiDb2Vq+gBRREheIe
GnmHzsYz4wIRcp4vObxjrzfUs1AOWfrWhML8jBEjdzsnmSOhEJAXgUhAqzEMcX56Efg7R/Y/MHIb
rMU75SbsxeibjK2CcWSz+8e2Teai/s2JXSe9gk+WYJ+BUPgbQ8kSQS3WAc5J91R/wDl2B2QpHoJb
iSmXdmqHqh97JyOwMhQo/4rdN6JCP2MU7WUY+NyBicggHkwLee7m3HDRQ+cVnX0LiGvbbMoHwP0a
AXkZOEgs0+5OS+676Pws/QNV2olboVRxlkB/WqgEARZW2BjSgzgX+/OP9zve4vs0yk+/HuByCdd4
biCplr1/FdMbjMVN0x0o+s7rqhPY5IT1DfPA5elmMoLQIWZ3KtasmVxS7yhjRXzOrEM2XaDNmzBu
JbLkwazlciBzwDvWv3Rj3rKODNKeDsYgj6ZXbeJoXhMUPRytNVzgP0ptuGSl7AEwvdY6AMdkXQlk
CHKuzsql47/PLG0C06Ar+UNl1Fa4wFDkyo70fIWCBCGBiBRkjdO2540KIWPh3g2vZuLrZo6Mkq7m
19MkdXPMGDWyJ5ctzZS0mv4Zv0pmI1a++e3SQ23DPgakSDZdhDOVr4c7cqEFJ6bEogETKR+X9qne
R3NEOgo2s9MDWh5IMiyajL583lNrkLcmhKxPY45q74TxmNAztJkcamPl2gcyXT4irKfpyX0+HCJq
I9NzRfc47iPc/remSLDQlVy9zqvK+Y3jiP4J4sL7VESJDMtq940/f3kwJK9pioA8HeOggzlYU+of
nIjB/C6t5tRUuUPmDJ0TZjftwggpF1aqcxNLELLQnW0HgJ5fdcv5MYLQpTkhEgBLa+NrhA9yryAg
3sb/wcTPAFNIuoqVASnwjZnWu/1mtvWVCct0zhnw3STyLIwZ7Z2fahY9eUFWnbHPzRPocDCiprgU
3crUACHOR169qPFIBpYD03x/dS3ZWvRl+9bUp+Bgz4vUEQ5CkUzHNEKWesGIQlBQxUCrOAsjJM5g
wy6hnogJsADEY4qdDn32xPs/8UlcXdkm3FGgzFCeMbBIrQ2lPtNU2q1OpoP5oUPPsx8ko9NzWW44
bEFiIZoeUBIRSfNv+SHszJILVGgjgNNXqGiqKzmLGoazEUgNLbIdm6If4f+whLxGVasaKbN1be0U
jf6OX6Vxao5Bf7p5wUWnRMfvDAqeY+syyMzuhYF9TezE6LtVSx2j4CS2ytRyWRt/93nM7/k6ZRFM
molB3w2Ubj8+lWdIcJePN+CeBIxzSsDy+fC6wudhu4DEmHagTtjm1oQ+SuMlWZ6yzlK7kCzYJs6h
QNZzFo0oSQXm7aM4w8kulLtPe1PbE6A7XpTYnRNlxEV4i6TFvaNZsrvs7ACiCSS+IjVPQZdKjmA5
XYUSsxTq1siwJuJOVIlMvON/lOtNZiuADRs/dx/4Qspmu4YIfQYX3bZ3PCfzdHXOOhct1mIGVrBA
5Fr0+xKsfFfeDq4u2gerN80Xgg6z0H1OcZRURymeOl26FB0PNHXxAdmCz47s52MhMUtA7s0A8tcH
xO5lTyzrQeMLriQdmbezkB/Y9+2lvvAZa7qMAjTNz74uBcPwRKiDqAi8MbQdyET0nBNkqBhf8f3a
2jdboQBVTZDRIA9P7UmYALun37ElF69wKY+RegspJmBDmPDeKGIETljTa/MW+zYfIXpN4hXkx/m6
8ieP+4tvQp5y4soA8B/0a+6Zs6/8OnUCJOwvN2dks3H03cPH/+QcjVYcAGoGA+qrTtmjGx624cwK
FvxAPTBinUGN0lbh74hN0N7VhTiGXLfoYtrEk2uqc/MrkB2YZj0pG4ZsYakhoXdFdA/Ky2VW95W0
AbB0XEIotfTJRqJ+D9ibp2eWU9TJTY9/kkflA8F6Xleu1dUKq56nqGAW3ezQChULb2EEqpO8rUjN
0mVk1ULrR9nRm1cyywac9xtJO5ipMF/eGrr/wPMcqX+nNuUZDkn1GagMs+4j5rnZ76N6AJR1ugJ0
xxpGcsNzD7Nk+1ZOX1tnNsDxS4AXkW0wXgyOshV7pGXTwB47COdH1fZ0ev4hXGI3ekSZTDYTIiA6
2pHYzRITnPdSfUglAC654NzBBDJFzhsmEWIQjw97uWTeqcnOyMcaw6KcaGi+QG2f/V0xlnBBfTDd
wnEY7EdBgquIR5fVFEMzGSR9YbjxeBqf05QfPtUQgLQ6UUA3gtTNwaaAr80r886jaA9azVC8Q5dT
r429NBX1s/+jF7WyqNX6RluEho9hfZzQMbS6grxn+0r1AM+sg3hbU0DjXFO3UWsx6Lv/2QyX+v3u
ITl6U72xw34i0IU62la9intBIoYU3E5+Y+by+Qxvo5m8yG+J6R5x2S9bRpyppW3DoWpBqXjILQpM
gDZzXxuUKbQN2eXFUbVDudn22hSk9BfV7RtvxpAUNLrnXnbMNooLX7r20S3IETMqPRMmoBYlkJ74
NAa+AY3NkclfbHy4Yd2H7vJXMFG81m1HPjHI1d1DLTzkXgHS8LCSheBk/KaHWTHaYjnas5ki9fEL
XkeLevGw/RxEgXb25bGZMausefYBE6qP2HR7Qe1v2oZiFZRzA1hK605mAwly1PlMolPDzis/SZiC
rnvZ87feS7ZomslrNWymGO8QMhS+QtZOjWFt+K90wMfn/7WYkCdhyaji6iHMwiravgxEPmKTCXMr
PkWpw6Rsyph+OYGz1Ri+Jf3i/57b8f3rCG/H7ZN6jwPp7SjiN6DJr58MGxVzig8t2SNjbOxp/zpm
2G0u1p3lv/nrNLXnB/SYrDl07LEb2Gw0WVAnSQUlrvBWM8uwF/JNNF1cTr/BGjx7xLrZL62jX8Rr
jWjOSlMf2bSna8ClVnJjZyinSzwEvWDFwsoZRYM15ZM+5fWbM/lgMCLW6P9bjy04e2riigL/OQ5P
G4KJFGCzXESmmJbEghtXkriZX6j40D4H+FPEAc/AMeD7n5jdfegruIkbv8Pt7w0JrFHs1wa4pkS7
kuU8EpfJB5ppQYhgZrqdEUoGWX6QYTM6drznpg6hpocKo/mn8gROE5yBYDfPKn5fjKsbOA9KCwBU
WNOWmPtFd3p7GcAMM5p8mPj8QxoLaN6cZ5EA9hxcVM0ZIZdFH7Ro3xgU9GF7U0n9lAGAx8EYSH+F
OZNXXn8kRzThVh+SLtxcqpiRDy46Rjuv49les9oJ5L6s0BH8r6ubIuTCFTycqHB5Ac9WwUBiKdUi
BNYn9UHqK3GCJrafWj8NVuqrRPJRR9cHSpQvxrZQySkmmYIK9h2HYc6GTzV4W16f1rNMxKMKPd9b
rkApCUyLcCEbF7Q3P5d9JLXG86iGjFCyiEIaAbHNgMHlEM7Aiddigqb4bL8Q5wIl8ZvCOjFKxtLA
gsr8W7tBa5y93DRFSGnfldMceKXjWRRChbH977zeDrGvHT+BpnLijw4cqzy/gwLzsJq+s7oMIOaU
/RFejBzk+UZcf2xJQD3x6ICNSuZ/dOnV1dmgDi1lCX8irAMldF8kDfeS35wSEUch2kq5a2uHwjUu
ubtupnICV8X/NtlRHtLpdsDmxrdN7eAT+SwFELjAOnJL3ual1v+dcKAwcNldjDPItbDEqDa3TvYT
65mkyh1AUtsDgt5TcsVCAl4EeBfiZIW7tkXHp/vzVKJCAQMFeStZWzYFeGur+jgxZomf6U9UTrsn
P04n5xJK73Mpm4CVhcCRQ0aNJolegDZPDTrriHvS949Oa3nR6zBK1wCrNm+UqU5ant5KvJZPsXXH
0nHWtKIvqaz5a49P+LQ74Gi3a5cK65mAzNRmnN7Isd1n0qH8HOP4HsbCxH5HsYC7ne8kzzTcks1o
6DdTlSrbwC5eKaC1YQTAjkJGQqtXDfAk9LRwwS+YhnJcX1wS1u11AHxal7f/Fn/vfve1lWvLcMQK
NW/hrI8njcr6vi/kRGg/IEUWrE3ubTim4j5Wv8SmNjzNAEpj5biIyOcm1AIP1s8q8QuivQvExjSm
XebszrzX/UrrfpQPTsAZrKFYWkpJSLFv4zl8uGLM3LCb3Roe3iWgtTSwP8f28t82TokR/2hNvpGn
RUoKBt+T60ll21NFuds27RvEe2/K+Kw2C7NKNK+ObGnza9nBLaYiDICIqnA4xcAm8QK/NiHJMtWJ
iamRBWDMF75h/kCvfY/0yimU3OoozJDtlXgPrZFO2/lgCrFsqOzOcumMJ389wZOD6xm0VnUDoOFm
m3oF+TLt/ZmXv02My6AmfKOrrwNXk/tvYtR8DxyV/Dzdswrmh08oVb++L/II4SOEqcgTOoFPsQnu
3qSDWL58jpK6je6LZ6oTKqNnwCFGTFHaGqnRFAjf8XlJ+uARYSkBNCp0Tq4edzjg9eRx0qTHMF0o
rggC8qkqLunatwr7T0ccuSVD7UrcgAxhz2PQHawcmcPnf4pHElTah91g7pcQ/Dp6wk+UDjnUHw02
muPutOWlPDzXrOLs/GjuHzokf8N9bqs0lhi5CV3WI0RJiW05j5ouwZLukyCjGKxwDVQkseLxkHn0
Cna6dRioweYAX5v/S2q4wYZA4kXzv1kSrPJhgv+hKQeA0DGxBLVRKXVt+VT3k3bO8yXYsW57iefB
RolbmJ5OpQHWYTRCVYf+LRQHlUIhFWJPqkS8byKAdCiDCDt4MJG9pYwtAzmxa7s+Gzv58cugUKiH
Ebq5VIr+Cq4G0DmS30jFTBb2zVIkfNMIKEhoK4C1kDhW52T4k5RVgGokkcUs2tIQW9xT4lTChCRD
If80tsS+rCZtxbuIebvUnohyTTviCKjylbpzVlVLYdC2KqUF0obFdXL6DKX5YQN3hn0iBazYQ8u6
eeBA+MwMelO8RLI8ZN/nXfUw6Hh7d8AXs34MeJ3KoKn4/HMErl8V04haEuWyF58BJxENx6SV2vy9
YD8fLb4TtakrKnMT94bzzVH08zqGMJ1m3s6CcgHBbqnqVH6mwfvpu60QrTTs8to2DE7JYoeSRBPi
DGI5eBQi9lTp8CEGIsf16zutbqezIdY8lVYwKHk0haygdrc+gEwpBmgnb4caBcEDEPRTXAjotnc3
StvKxUIrPIKTisV8aZ/Gd37TRV0/BGFz4WBctBIWcA+fGv0trZnSvSLa7JHXo8e2KLmjzEhdW5/h
UYL13q0gJTMTVrZ27JgZva/gJrPAWmVIVRZqdEvcr3RmyQD56bRrAGGu1uZlTPQ+ZNbVD7+9cDaA
y0sVanooe1SXB7DNYzA/cW1sk1QMFXOA+y3cgSEEwC8huB6t+cF6wedubaGg0e4jeO9IEeE6sZEd
ZtjtQniZP2nE9DMiyVVRWa3UtiECDFx8/Epsk9t500rKkFUj2D7u+1sTlj/V+G2jw3JO9mql9lcD
L6VvOmzTTCpMP8Xt5xQkf98BgognuJRxU3hFZ8eDa3LcKIvnFx4073IFwXkexATN6ksjPX3kXiLG
90UkvjJSqaZMtExNTlSBw6noEd07oEDJjNzmqxo1iXbOBEvs67kQ6TkfX5OAAosuf0enGNWL9DYq
cno5W4neuvO9xuzqSwid5mxysaVAoUbfZeW9CXIOWMXXeyTdErCuD8G69VUOAhJK0NjcY5iXOKqT
lkM2WUBRCpeCTqBlyWr6nL8fqBW2BkRKiF28JPMbJRikMq6+y95pCsWvVbOl91h1ZweskgvmDIO3
folEWIMEUGqXY7K25zd1l9eC2JuJ1fQmOiOmHqVWMMMt8jzTn2Xk1a2KxuwSZpFtgvIcqQ8dghsW
nS27Ecc2fsLrlFE+RVeRuAj+A3E/KBrhzIsCPsAe1azV3WnH+1latOzWmOsl1yVLcsu/4O7i3ryX
Dwa06dZHi4S4pcMUpLp59ud+sxaJL5Vnozl/6eZL42gT1U9zluDpQ1pkMZdE2OOTBi6mSh0oijUB
x6c06tcGVtw4IA1FYcp6/j0O5p8U5aIJ87zyvBud4/iltNHYvzkbQHTSkw9ocQYonEvKcoivWciP
SqNF6HMqOA5vWPFAzL2R4TIKq3ZsJEM1zm/jZHxGj9WlbkJ09Dot+lZowk3/Odett3kXk820vwlk
gkXe02egmJILUJCWBSLxCNSDLbNZSn1tcyXLT3AgnKkb0PqTtzJgKZTbRIcbcVyDCGQgUDib5OMo
YrjAdve3eu0upVy8Hy/7GcPBstMPIGrb4zW10zr9AnAqudCfIbrRMTshk33Bw2s81iDlYh/nOvWy
p/Lj92MLyJRNi+YzvpHbutYXD7UNjbZXdTv5hbrXkbXp3e0MArS3kSGST8gQdj4DapKvsRPEF7En
MsHNmqzqHFwA5cHOEmwnSJJ4BFAfgLRBkyuJO5LMnRnOt0XoXhjCqwl/1DkzqGKyrA3bMFoGOkmg
rL7MMsIvY7f8jduYf6otYay2d4MmKU6XOCDlMC1Hsue4M2HGUI7c8AEmI2ToavUJ79eMRcBWpP9N
VZ6rzPrtRydh16dBJnpoJyzhN7zdqzNgOPujzhjcnHlnI5lnDV3B75qOhN8eYuj5xUrTB6vcFfQb
ICRiT23inVUakwokq0SCZQsbgF20i5wfUed4eYFQF0sasX5uQRCtNZ9RMgxuh9AeXNBZQyeugBmu
rEvBjFGyn1INj5uFVpT7k/ZeYVdxcEGIPFnDn+8n/Boz8HIsdo5epOSCbux85c6hBpC6njK2Zcqm
tQDYc/TXdo07apGOerd7OCQSZm7M5M0LI1zbOR70pFSqKbrTCO6MC6qbesaoPeX2JQk37W4B2Oik
ZuKQoQ3wOINjeTEkaqIwXtrgUsOuP/jBoLQVhWmcx9u4balnsRQa5yS3wDTJl+7l9Y4hWM/U7JbC
wbguDMKnkxf+ktJ2AnzQ3RaXSpvrgFfh7s2+nLW1e5tnp+KUPICs9ynNf7Bah+Ch388yjMKpkkdH
3N5gWCLSbOV9w03Lgw1Qh4zJtT53KdRFTQY9m0Wgc8IUoSCMMDmrr5GdhisVYBfG+OZy/gyVSAGX
H1W9tV6qcD737SJV9l1eAaybA8n+TbdXhQMmVCWvqxbd3eBFPczX09+d4H+B25SADk+LYG/lkddu
vdtbEtTze/IRANSo2ZI2o3qi3ygCDbYBmubVuq73Qgi+eRADzeOKWrr5SI1OsCuje7VbeCM78ULK
Mcg8vvOtROQiLResGhjs8e0zmJJa7GFLGuridAV8MeQyx77PQuMUnnRDLdKHeywT+ueINVj2gezu
dva3Bh5y5VNGAl7BWyuHAz7Ak804UAfg5+xup0TjFyXSukjWaXjx6poZZtDZ0TBFycLtvbdJuPdE
Pye0MwAPwzPew+I10+TfH7rq/HkkN1BNeaX8ZwG/RexDEZePU61c3Vwt2nbILJQIPch90mBrQQsY
qiKdhGzT4467Wy+/ie8B9oc2QTmKdrqcHlqbf9HO5iLooziqSIBpdpodbXPbixEg71I/TC17zEnJ
SLwYSrup8yrTlciLelFN/bnSsce5G0sK/rE9Ch0DubVSVr3fEwKuwJ/uH8v74kbVg8PY4Jy/reKG
DBFHy6412AWsvCdJUK882U20zllMTQzTnOSMjuM45ye9ukStRWOnwnaQ9dliJ576uW37p79mQdg3
hZJkXUKFXljs9NJRocA5Qt3bS8JyMbmOGQVvVdYEKuehS4Wwnq5PBzl6XZFM7ZvVc14Jr4fLS0qL
c1WHOfM27T1PKWx8TgapKdemgLr6a3dgjj6JKxH8OT4phMRdtZEDn62QGnJBkkf1h3/zM6OHZ6U6
D7MNnRyFR+I0OpRzVplPybsHMrEu1vmMvSH7DMsHnZJYTLMeNTWxPvITgyLnbFHOjBB1tLVvlnFO
psA8Krm+K61pY19Cu8mdoyjNpzIZrPMw/0tgiTJdmfQH7GKlLWQ5zk2qycxKjkHwVlEVglzl0UA/
3Poxb5qfB5uqAfTT9xUuXTchgNjnkVA3wBlRIK2OyODeMiqtpxJ3GSYXfcmXor2mD1Oe5BrmGG2v
76OaLbxLrOa7q21quW6/ydkkE5m0gVkraTT5tEhDqAVwRagNo0yg/FtiilzouHkSel7po3AV/JQp
eno+EoRUS2EGC+xGrYGPF3ml/kGtpebA3ICJ1UDNgYQ6LldR9nM3UjPIgWjs9QiuJGY4tr7WoQAL
jdLvMEdpjpAOStT3xaZHkYuTnffF22fm0E3BZuAXUFNMqdXTnpFntwhvopYRUynCIr0HUPPycNul
27bNy4HzhJOvI438aDBQXLT5SGSTtTFFEaOZCifsItl9hPELUKiV33HFv1X46Qw7FtSZPLYUKC7c
7R4MjSKXBXtcZFUrd9T1tQ1OjK8vZuQ1pbO1Uh7hLdY+V3xIVeNDILBxSRW9fI/P6Ek8tvRtxxSK
L7Q7CBOI4ypX1Eh/3syQNACCXq7CM3raxI38JEaQiWZU3uHC8rfrWAlxy0kBHDaxI0YvbT8xezTU
2qQJbEpbsfqr/jxpQZ0xtuhGNe2TYjWp799J/JbEqCP88MSsy1mI7fA9RYa5qCoDz0Rrbw8IjFvu
Yw+qudjiRhQStEXRsEEIKOXITGSlqzDg+WqGK1yjJ2Y7bBMT+z2OBkPsUBmuPsObyqeJ+gHY51N+
xuyHxRP/KA5OnTCf6j9WvdYPbx+63M+eUxAuZT9IrNN5e5OfZZPghlQJ0DUsPpnxk6AVF1ux+qGW
BHdoWxTxZobqnLQvkHoyIFnoD8JDNP8t5VyUr7Ceq/RcsW3S15K0FrphTmdH2+eDd9Le9fh0KUXS
S7pf3HM2GCNVvFJRKfDj3rgBVHUddyd7BVPATeZCHUU4ndU2fSsGEUK/e+1xdUlOqm0zkg98vkqm
unBpE2ZPd3F2H++ahs+KtcnBBigWDn3bcoDOksa3EXnbZEz+ypDD0gux3GtpiR7Pq49HMXxtCKvu
PHk1awwkB/jOOBh69jgZllaBLKwwwJy8SfB+KKMtsa/VulXK5faA21JKMYUyxlWM7gdnrCCsVQ4d
4BXzzkmDEOlF6FjhRJUn6HAFuNgA2/2WPZ8ynf98pn9gxCYt3Y1TWgEtsAqT4ka2xOTsvxhOLypN
zKEl3oeUOhUH9zAyCO+wRSLATNU3Nf6pWa0NQlCW9BqxoEHzUUYy9D/ojc1jpOvdfO79o6AP2KRF
KzpZ3Opuk8JlrkAjnS9gnYj5/M12MHbEt4Y0g66ZDSkWfIVa+/HZpN8uuH+LGe4MFrCeTbq2eunf
sh1OgPhnD/Rm0nX0MQq3cD0n8QegPK7hWXvRYaZTqBS1FuHgsHUbjf3ZLA8PTw+DNVG2ipSmUdJo
q3SwbZFQ1bIpq+VNps72qIdLGfNPPpSjAQywf7tYVsf5TwP9hmwxQLK1KbSt+QzN2WobCrSckS9D
kVcuZIDyVHO45lSXx+hEGF6kAGmE0clIG0lsHBiWIOM9pSkyeTkfE0tSBdJjFEDlvkDcOPnlzOzl
v2BcmufLs8qZ2+K4P/JO3cFYjHuTejz0ojLtuFm/yTlfIJePaFlP6tNhZickGhyWIaDN3n0Po3f4
rmiauCygwOereEbetqBVNuaLxLVhFx9Crtt+Vqnoh03xAsBGq0gW+4Qpk8SHl9KlQnyA6B3tA5vx
m8SEoxnZEgTDf9YZEnC+/W+3HC4mweJNeXZMV7MR2dpLPoQncY4uO0tFKtx1GACG/9AK7b22eBPX
QXUX2o5yaAf4jQaHmtsU1hjMCfq1yevsChwW12K60RZSVQQMoy24k0YQ6KfMQAWfwy9S/OYfRWd0
Izb4AjXxymviL8uEuaepTz7X7dRO9S0y9/EbgJh9w/Iw2sE1M94ssUKWb7J2PW1sIQho528lUkfd
Fu+rdbFzlivxvHGR0XjgQ3WyTot92sx3h8SHznj+jeSkTZAdrGOLgdF9blQYRTES0T2ESrdj9vaC
wZzm3Phne3NHB/PG2K0XzxwT8dDtk4EqqS+9LEgS49tI2fZGXCUD+YBfoDOG5nShg/l+PP4cqoC1
DW9O8GhJTLCnb8jpRJ6rRoCT4QywDlGV31cMSYGmabw9uvcAMSI6xupWE/bG8JZ6mbwLbol9KKGR
LzNMi1ACVw9LLeABGdZDn0wHaKZjkabliCEmDrNiB10m710BT0WxG0FoXW9qTZRcJ4rMSv7w5BRX
BGF6wUP5ZhAo/DMdzQNXbM7EfNS8YrHafrT0LAGXJ7s2DmSPsRQmTj6GGwSnh8/YPHdLRNHqbH14
kL4VTfYypmJTLrA92cmIbGkTkGB2vDx3hVCYL2yyBX1ggl4BaYhnv7iVZ568u5danQRpJj8d96tI
IVQH/fViWxIIUedequUyEhJttUwpt7bJmvkL7OJNPtHgalZIwTcNqouB2aAR4AiRUfkQ9xIaHWoZ
LrpWG+M79SCpuV2NUqq/uR/JaIy/0ZpY9pUq3VjnXG27x2l82Wt65pbczLoASGlJA84p107kEIS6
4QuNC6L8hHrd8aZavTnxlkbYCso+aGARK5olqe4qj7oOc3l29tbCl32v6/CG8wJQFMzkDmvtk2KP
cgkvL28PccX+I/8jGEe9j2l1OclboeRlV9Y1kUzMSIXQX5OU5TSDiRW0mD/TMiGFhfgDmIFe6mb5
SLEUMc6Hx9c9ISQCfxl2UI7yXMKsjHFSedMPr7ncAThQOQV+KO6OWSLrZgJbALqrJEbFfbuMHg6D
jSCHGL28llcbvOB+di6UQ9jE7a0aYVFjneDfitjh92otEA97eJHs39utxyG8nT2CXRkS9eQPp28n
N06cINkZU/A1WgPYmOLRBoaWxZKtrew28MzBN72CTv2rt/QX6umzN1T2a6MPfKHw5VSZA55TCq0L
eLoON8Wn2dzxZJKSc8MYZZZ1GcN+ImJcPkuuEaGArhb2yqG8umg5wdyGM4uqr7dCOeoiEFh1At7C
2zzGP+RP73mJbWRmdakYpUulFYqk310IiYbab5OR3CGXC2/9XAfKjYm6rQEyz4ZASJSpx1mIOn38
WunuzwnoJErbshuhDz47sD1DQoSZX2W/AFh+jayWdd2PIfG47dWhVv4/uAI4NDjgE/jP481tmnbG
Sh4P6CCQckXjDeRKzsQKOIkW5Y4bzHOOzoiGrAMyTzem09uXfpF8op+p5KqTCRFmc0/OO90YRB3h
1RIX0JEplcyWLch2DOL/yOpgJFpDRKGoCrNeRqsgWRiZlHEXQi51app/h/Wb3DBvuk7iXI0Gzwq5
Dp4emhSubJeW8vdcdHE7K6mRIeHI0CWXW3hkPo+LSiMjCYsGZyDf+yWaEwHWq+1u51A1acMkkc6o
xgloco7/POl2k9Dn4SAj8NTLCUB3ltuMZUppqefpQAp/of05zl8pqzICu5RiH6AQKs934Ay3w8RH
qcdhAcuUrNvti/xbhaeyCF3B8K1MvKH/Zv2Z3IK/k5d1aZt0met8owkwPAMXWEBvv/OU+br+zhpe
k3wBS/pnaI0ev7kSQgvJ/QyTluqo0fEk6hli6/xPcJKHZuu+cEWXdV2kkHnWk/7aorLfZOodxUyD
L8n6GVNQKvPcNRa/HY4q9/xL0yKlxU1Hz3IEFpeL0ULLrFbbWsIDNmw8zq2FYCCj5EizGFz74LTC
ll2vvE0E1NViH3R3j3HgwRLZfSaqbwoGWEJJUtsHedF5GiVqTcbbOjKQIPMforB/Qcr/lPOeamT5
EozAfrbgNu0PGVinPz6WOjkLbfUSdSLwbpqHOyHEiWLosRsVwtlVYRWmu/kQIUzRUssMFv48CxZC
yETtW1ynpjbkgLonau0Ib+M+0kpFlCxV36ixqF7EPkmJyKnY5H7TfW560KaHTxBWWIHXzrLwV7xW
NkHQYiwfSbIci/m9a+51WQ/aGo25xL+sObBKKHrbKoe4ubDAfurmj0Oz5rzuqTzN+Ytm/XUhMScl
Nd8hRsTW3tgSNjxZGeswj/9xVLHVEEMAJ3Vo4O49HLe3x6rUu7SXb6CDmf4pCK3GwTnjcy1jMhIe
BHcv6BGzff3U3gPcmozeS4usGMke86Cu4Ova4Me8INISPu0ZAqzvhlahqFwjsrsEhg9JUEAWeckm
42bz9ARYySzafW6SduwjliJ1KLYNgJOr3QU8oCGAxLEJXDPdJqqsixZXRNvsVw0dfp9W3rXRh2a7
ue2zNhxv2OrhPXdyiziVoqX5F5Q1eGRaSXPdF6xDbgUNf5MhjJVuWr+8NQSe/j/JSuEKjYhnsJpD
+orNdec8ziRqI+65S+EWec6VSnWJJWBoJRzYy6YQ38eP+BuCS4cX8Dac6bBCXuUJb86AdEgFE3nz
Q3cLhvtk2WR1i3Yk0FPI/VnPTMPuHBT4rsBvFGzCZ8ATiPl8RAt0rCXFfWPr6Pu2gX3s7jNDvoaa
IGdFkbjkRpYBD5ARppUEyomG9SehAEuLg16OHZmz//OIV1VXpOSVFmCOr99iuOi5Gl0aU2GPKrES
VbVSEbQetJcSUs/8FVhwL2Dj88vr0Q2rGf4xvBy3rwuY5o8xg2VWVlv2cgvzsPWEr72crbyMZ2S7
BB3DDrCEcNxINCi5sd2XWmGaBq+5Nz/uXYVvcpfH02sCZ0tcfXVKjtSg2yp2AXPme6CtMiP5VoCJ
ncaa1VLA2tHiHQuyYzVcDOLLRml/5VhgPdUgRbyw/F/EFdmnyiboI6nZkbQoDXffT0HJf9ZxTAQ6
1J1D5xDISk8ggksB7D9Qekn/TNEUTr+UHWUWWMGnx1pYJZeuecLWIhUxM5/YcmvzsioBsk54l8UR
9kTKthYhDaGDt5hlug0nVpVVEVj8FSUSessNQIMTF+8SqX5cpScifbLaLwzjm9o/dWnpVN6Ndbyh
oOb1tvQ6xeiTt0wJLzrLLohOEEL7GjVcFoIaVHuv6++Uf6Oxv0PBmnmopaRIcj2zTgdTervkeKE0
/diLPCZSp0bBOHbgbLNK5e6Zeliy5z/8TEnPtGf9RjFtZQ/0IKgKoXm2ecIA4MQCb7cXJ2qV+jFn
bRJnfUlEFkxerBsOH/Dv9Hr73bY5l8XbCsuAL5FCwRlckkvBjdsGZlUyUmb68y6wy4UWqu1OpSsQ
zjYOnpXDHuzI2C31yTGQuBf18ifN6x1pTpiCOJ8ZjJavaFzG/2TswuDyaklymGm2JBEoYTx+dYrM
pmAADD5pUlgxzTPsZdanTMG6xDRZkahvOgcS5Djf8S4fjSQHX7z5z1zmcHhIvktN2zdmK9ni0IlF
CH669dbxD7gz+EQnTOghtsgNeSFcvxpvuterHilMsMlHqTuJ32Nq/4U3hbbhwJT2VHQtMH6slZJb
+dAg0Fo/rGHJUMXeIEUIetprDlVQcN5v6weKCy4Kg/5PTGQnjbC5+m3cFmhDCnfkKULFhj3BPF+4
wvhm9vKSYCsKUSRr2z5X5KJXyjffwDC+rV88cP6rPBEMSgpQkGWWZqIoagfGn9vI9DAywvx+9lIN
w09TTnM3WjnWJcPpQGhjfE20fUkH17DTMU+oTGunUMdFHw4m4KzdOm9kymxvDWpSsgOb7evtR2j/
NydxjxjSGqNtCGLeoctMcVkNDCUw/V7CEsfR+UT59d+UeeM45ctCOec6OpGEBcKoTa2+W3QG60Go
f5+Ys2/DlHQRxAw83dAqTAlZq2nxXzPBWqf/2hTWYQD0RmkgM3hN5M5LX+0DbUOK9h92m9P6gXB0
h+E8iWdngiYfMtYFB6qt51UfQl4QeXUaaab3QvHSoXWrJXgfT1jxbZWfCyRSbKWkBB82bZW3lcuQ
oMzVPwzypDRsLcnkGDvGcE3upGDhdleJ47bZD1DUzVeoy088sHF4/L9g3S9H/cjSp8o9EobvZBh6
HU6gX7MENrgLt0yXx9+VXbPxjgGdnae2f6N/cCfeCXbn2Le7rEIEezXBnnLsBoVYe8bqtzxrCapX
lkXy2CMs4uKfuzanYn7VErYUQgXTP1NowV0KRE8wTAPB7Eo6SVXM9BdlwbOO925bA831fu8kDZMK
yBAZB33zMJdIP05V5DO3u1ZaiVb0ixmOzbE9jt9U4OMpneipcR/jCreng0ubV1nFmFv9iOi1dZ47
swyn/fiwy669dsoZKBgsjHfipT20kSEMMRlZwukwY2q0uc6sMnIrktrEZmPye/yxgXWFtRmrRiRC
7WiPd/n+Vf+Yexzlwmy2AHs/QW4uKRzamODUhuvAn0pH8fiaCMJiT0qUnEUBZHrJfa2dFNkq992A
RPutPcHceZcM78EaawCvvW7ceRNyVHDgDMKbvxUuxrkQH9q1k7hvylm7ztk7vrOGe50v9gspvVkN
JnX3RXV/m7MsKyY6I8PBQIP938WRdfk55i2/cfyFaP5vWd2erA4sHPG2mmKPOoWIiuK7SNdFSea9
UmmYFoN6tCOnXYQe8nsjVtm8g7LlT7nV8bk8FAts/NDjOajGZoeAacwN74QBZYd9dLSVpza5H6Dg
5AHI6YBxMsQkaMolX1Fue6hYi+5R4vqIeM/UavQ8KY+iD8m0dnt13cJhQbQPqEWVpxRtH5ImNxIT
s93mmHGO5o7KOr5RACOgzKXz5uGWE4AJDPZwCLyw9HWTJf/NZ3VTaHoNdr/UV6pR5gYGqz2bt5CV
xj5tJq6SD1kZyFarnEYV4IaNWaaIOxQDp/9nbtC70C3m4LOiokp5l2I5LDB7gz/Gxk1jSVPYwrQ4
HrwnHmb5bGaTmQ3G5fjdFKuNqHfDUBmkeEXxLNbDB2fJa5udzrvT9omPF3bn0oJfD12Z+6x37qe9
IW0V10Y39+GiypRJXDwd9q4iTM/vb7YJGjggdUuTDkluJ0vyQB+5UZFWnNNS0883tWPGVZZ8Oy4S
4fO/+OgHi4PiOiACP5hEkEcdjZpygfoRbXLVLoJj5X6t1bOQf1u4DoVCKJCmmXKbbesBB34ijtda
HzAf02c3C0Yt045PkscdzFmPIQcjYlafcOllJK6sDxU2znOmidhm4NfMwBjn7/UZsBUQ5kKNUXP5
ANmJKFpZDLmF8pRlLcam/e9Uu8E6DDVfiHzS7Ci+uhEBoSJDUjaKGmb1I2TZ9tdmnuHnkKHGHWeS
Setn9PxKDUeNDpN+97wJRueDXFodExe/ruXBgdXoGrfqjfp9+NYmFbwSppgUASKKrzSNjtrn0ajR
v8JymTKQ05wV6CcmMwSCshwhYcxMADaV20AvSivrBQgyn5IdPiEw6yI/ARUSGJXUVspPg0JtyZAe
E/UY+aeM05YE9pIwRcT4qs/RNxPr8ocPMaPMFYPchRaN7yvfu3mzlFwd+lN+mwNWprOWlfehFOtD
dbPrgPGT7RYuwdTl4AKZ63SxPlrMTRCzgHGic9AxcRDTiby4kdxcFJwqu+dvJE1aErKHe1+Uj+0x
qchblOKhIVbqLXmWFliCUdVqSn84EigGFA7GeZlnzgm9zYq/V4nNqoI9Fm6xaUAM9Gi+zjhwxoLy
7337rLjOmOGlDFEN8hg5iuUSW1Pq0jM3dQt2T47/scBBYHqo4VsLxikNuZYHOSXrkwWXc3xu8aO2
MweaL7vCpLdmdRzbYdZhKmXt1uSdTdb48JvbylSoAS0lRPcRbWi+50oWjW0LV3f8mlNSbc4ZnsI0
lZKD9PDziV9wFZhU5ZkWTIh3RXFcvcUktxtfvUEfufqrSTdWR0OJuqFxzArwWOh421AxrI6bChBF
o9g8RdA+ryED/ZxrRh20YpoWtcFTqzZ/vzWedrqzB8Wy+7AgCNsFKW7CiFQOkhIbIAm43rdoUtlT
DGFACIi2ghpnKYDrv13UHOa1igxZDc/quzKcuiXurhQQLIjWqhDyO+IJ8j71I9+IyFM+Z5zEzTDS
Q8jIWDewQ8DytRbGH8mdnpa+0aUqKDtG0wMsOnxBj8V7Ec3LAvJT4iGEUc9qRbh8m0jcZphKNfwU
8vNUG8EdSA/xveJHbWqs58o6k/fnXrUVrJ2nApUtYNsYxHxMUQsnmP7xpJESRx1dga0cc0zCQXx3
AMzBJR6wvIYuF7ZO/X3+UBHUv6BVTjAGWnZudEuD97PmcnQzySp2WWZN/+m6KYUU7Zj3YUDEN4PH
689AJP2m9HawRnaaC5cavp2XdPUxDq/PsjU9m2Ibq+DcAV9EFhNGBEpeWFmWU4eiV23PrUCnoK+o
aD4+MJuHdvbvH6ShTEsTX8Pc3b2cdOMzNngKXI9sqPvqGfZlLSpSbgx/dHPFRB26buto0MKesgLg
uNNwfJmjNgtXsX4qS3myCpY2y3Bcur99IONHmzOIBtM3sUZ9ep6VlJyFry8xbhl0rs4hYROjWri+
2N4H+jLRCuzENM+KNdScgjKq32LgHLi7aExbP6janpZFAepWk40EKy4t/zxPrWHaQ3OgLf8iPE3U
rZ47J5+/E+naJIptGv6of50s1Xnh78ioCgHr/rWGO7kB1+r6Ua/ddxrNr7fk7QtKo/lq0sk9af5k
JFWsa+HgZRf/UytxBV+EngaQvNi1LRiIAsAWelMCh9ESU9Vs3hwQ0QOMP7XgnT4S4EWpr/I1huOQ
GXkvbsvcsYKvuEOtml5kibp2Mtb1Cd8GWEzlHo9y++MaZhc2PWOobQV8jTB1nWG5r3BEOeVSxreY
176RpOAr3mr8eUhzE85fJENeBdUQf6RtRX1Ked88u+G4coJdSLKgep/yoB5nMTfCLWphnqd3Rq7h
mI6hZq3jsa+eRaJNmALydHOuKy7C+rdsCEWCsmZs/fOR8eAm9RyHjaZK7l8F/weegjLWWCeyczQP
S8G7Ee5c0mhryTG4x69q15oD5zVNZMQ/UT32KpYuXOfOlBHYRPv59dGcyF2OlWIgq2WAJyCunw1G
tiDfdnEk2hesQ11F0POeFxYrUywC21q6Pp3sDGQFUjSygt7pws68npJtBPLI4HADR1PdpQFqg+9Y
zwHikMccb1UJv+giWW9TSr3isWbLiseRxB/o/0H9CEU1y4kMtMvD4mle3qcuX1e/VAaF/xDjqyBJ
ynDu0BUG8U+S5D2xIlo0wal1GCJ7PNAPDXTV+6QjN/dvxwnZktbzi6NC6Mu7enncxD9BrWIin+II
m/B51Vnz9Y83qBh8teTWyVbHSQpOs18fhLagR2X7PU7DkA13feNUJ6r6F2DLRPfhPvhkkoNpi2Cc
f7iJvckVJDT6sG0gQDpZ9tcmqiLckZLUod+vJdiC8vrpK79gpTsiqgqc8DLpntC4wmbY427TS7Ys
1WFRSYvdCcU0TcmMZwvDF+tbeK1/k5fK9VPAXAbUEG5JYz+pIqBLggwa+6OLhfV3Z+X1t5/jX74+
SZ7PWEaonaUsuXW4kfa+i6TBl5RLJDltaW6KHTNK5vv3pTTou/zu5Q5vLXoU0YnszqqoxxSWLQ4s
cIkvwzMpEAzY3/9+L5Rpu2uiiBiN2VN77MxjVRszONBD1bFMQMPitw16oN5axNYaytDoXO1BsQOo
X1sUQYu4E0BbNuVb3j+rY5uylyk0g750EtpWdB9j8g+o5xNo8vOgeX2GePxCJeRwfCVV9R3AsbZA
0hEfJmPup8V4UOIy6JN0r10AS4QJdy+LoIQvndL19iyBoCyOxsdyYezMb+1Jo9aRYiIKzJktQWOQ
sZb1fTL+vKMQeb3kJ25aTxLoi14wJqE7d1BBGb05oyW3BeBt9kG1NwDJ37YAde3hHfQcb4ZuRmut
j764oM1h1EfeNFBJwEooTP1orOaR7dXVrhSowSRfRhT9RNhmeOcYLTTVZ8nimVGHka0AmVHauiNu
+iH6cPEQKAPF5TR0qX/4vU+ZkA/qXzFT+qZcYYjc3X7TgThgdHAKL1+5L8NwMnx442CZ/pTkhBB8
74tZsSYh/febDakdaPrucmEzXLUPq+tVtW/KEbGr9Jo27KVdjczFpCs+ovV1IEP87bKW6fDzvpaS
9j0Dn/egcfsQGq5zQqdJ1desreCOYfUB00RdrWMDbtPDQ0P8OKavEWdCMs+o7V3YFkC8tR/U89af
yr47dLUkt+AtFvp0lHMBUkfINOlXEFSxlDdtDuNCBFvGOAhXE+5+pEtMuxSaQa6Q5qMrSq/5hmuI
YAnxVNYgqg0IzQvs5mTVcIC6HLg+6lYs1BVIi3o3iCDOu9lqejQZHbdSlfcFDzwsL5C3iAtTnS87
G6VA2Dha3kRwl+z3Q5MaFy86uXih6zAUax7dMpu9d1SwvNiENsvezWqPZqy+9BLhtZ3ND9Iz/Vu9
t1YPJAGQapgdzoy8fENFJ7d2QmoP5kbFK0jbN1pZe/lWWtCBIhRTupcvguQzqPdsdR0ttl2nO6tW
TEFxelBHkVRabOtnpiXfGEWM2CUOht/t5SVIsvFj8M900EgNYmDlokaey4jsSg/W047M3Bty9ztT
Xx4dCIrIVIRAQYJQhqgGyYNRbWFkoVB0UqLp2/ByA/zzhoMgH4/S7jK7xa1oOaqmHunwTSv79zEQ
4iMaKkfQeLlTMrQMPfidrdsb0Zd5wns2vxbqTYW4pdp8mR8kwU/GWj8lD7AI8hvJ5luk+tgkMu73
aZKVkfR1mqKBwM9nbqJezca3QbJjrsirIAwAqdjffeEH5O3SQz23TcnZ8asI7u8hDh9P8HPL3pTI
3m3y0gxZsXBrEXkgOMNqLueGFvMFwHVxYSVqKOYejiF4YqdmOkT+O2fWxAgKEUtrYJHFRHcEPQLG
0EqFpbQ5tuA31EXw2cOllZ2V6/ogij4uBATwrsl0SiGhnU3Tph2hidPd6aMeNmJ7qJUbCRNNNkFq
0n/JCHA6KNn0cBVODPahLg+wrWZxCpeUzrSUG1nXWoIAOA2MxFq/XmxGtBlEWnZ+wgVZtGEUpkzG
h6yBjJJIoxL8uVC5ozfbAUKYTdqqRSsT8Cr8nRpvdDONl9mKTzu6JT6BzgP9PETi0S5WVLltwrdd
zSDJSKuvL4tuox9N25IirKuP6hTmQi892jUdCZoX89sH8+7gW5bRK0tMPlckkzSN6DqZRjGFEj32
3Cy29ZXqOwPzOtuPMgTQ8rwxByKVLbhlOqC75xTf34fIpGSRaaTZJNtibvfeQ7eaSKnMVY9nAqbO
lPVKSn2pYL8VKpdKS2Nis9PraaKTW4HXV5gvvghSTNiwhR09XvdBNlqF9YCVLi+nsd4VCHviqGXb
AXLThnSm27Rvr84udFuayebXUaNPVmbRjOUvKhKggU3l/FJKejbpQ5li0rh97QUetkUHgc2rU/ug
cGsGQKvKqBfOQ7v9Wvjcn16FLWOSwaWTNQBInrkLksEwqBZi8Bh3aUKyFYhfU0qGdLGwNI0cmE7G
svDQfg9CKx1T1SdddqKauYwe2nLhlwSCdY1j2uJv3M3/rlm19N6XA+xT563+IGweA2ktkUFAiAtt
zQvmhvVtVwzZjBVmrssDdLuqwA5p0ewSprDWv30M89J9Koz6nh08fKeNJo7YYGWn0CwH3+EJuy19
ZLYWui7qbkLuEvi6TS67ItoIDDQrBGygGD+lF4kwtBR97Hz583uxUgRG+yof3FNlFAhckDfWfNOf
8RQ0PHRCFQ2CA2X3zofABHPXxQ6HzSNdarMKWdWVr5iJPgehqOe1rIm+hBk2dMSZXtC8NsY8A2lz
aM8thdO4dOVWgDPP5Ecn73hO8424JEci64ow+PN+Tp2KlQjw6tgYYWp0i4+DXBvgVTnVRHXvQAw7
FXOzxr8LzLHDT0wxSvnXHB0jLc8RzsAhWpuYFHv/x/E7iCbCFs/wwttBLEBgjR671dHj7onY15sX
Lm9vFRTL/AMfP848s8dx7zG5ZjQb8SuBli/8GG7vAQ43eeUMmMl493FVWS0vsuWLcC/AhVu/OzY2
XPquBgGX9so/792+RzguKmhCrt/RWALbbCeH6alVMzgc9F1L/XxszcNAT3yAuCKTGg8/q+utM/Dt
PP7k3y21McKYdjCPM+XDID+Ib796ENrJc5wei9OINPzELL3D6Y8kDmWA+LjLEbxX2o7K58SnxeKn
J78WkkmIf+RHFi+g/D4pzxPy7fygRIHUQLBrdTcX4xvfIeXQLLhn6q73AWnb3vjClaKwkUV2jwZ0
bGgN/DjQSOJB/6uzCAZqeWI2NF4swH+YAePFAb05X9Qw4Q3M/MUOB01JEAdvilNMosWpngMxfDU2
6ZovvKPc4sMwksxjOw1mPTzh9bf8dp2aof9WLJmpLqLVcyKZjQykOYo7jpX6OChczjXMsFAVvFqd
KOC2GxXc5+bgKyG0+NJXBNGr1Awf+0r8kDYt4FE3tqg/gihHsCS+Rkr7n1/1vkz8XoSQ3YCrqEtx
q+bP/QX2lYbWKQyuMKYuJXlnyNNb8G4BDBxmd+fOAh3vvHPIFWZeLDNy2fbhXI3FoAgbnNb3B2P6
5zS6qMeJ6j/DJmemoi1Ym5IYIKC8NxugKViXEvDzSWxd3uvFU82hrKiMrYlvwwTbBtok9+RGNlgi
yVe5+sNe57AkFTPRnE2WEYJCh7KrtSz7qztW3ann4FR0wiglSaKwxx+z/QvqY+M3hXp8MNbk0Yly
0fkK+68z5c7pRQ5SzHXBGPiX8g7ZBr+tERZknoLG1/Hdo2j85TV7kHSOY72WVm+fYVhal6SRQ6p+
mol4vRCXxkoGwmDCihBBq/MOPhOgxKqeoE9GlrjsXNs38BOiU9U4OP0NeEm8eCcNuAT8c9O4W5vt
3E01noxEKrK0g2tVhav2fVutbQq+wq6Clz4+FH3USR2SATpnKSfoX5aRe23cmpulwR5hf47C+qkG
Yhaa3FHaROIzv3ZtO5gj4FXXK0+S8f0lk8pYRDafSOYaIu2U5Fzob5NqalU2fQ4+U78rCxql+ORW
ok4izmGVm7K6H2IY5YyNp0sKsMYPk8P4kWgyj7kQNUnscsFft1jfJN3U4uNqiiSOBRmAZeSK+1mA
G06qJ8VGO5PI99nt4fWCrosn3OhaN8Ah3ELCB/I8sJB6EispwfHqob7w35aQWqd7M8QjYW5Tsi+s
nhtsH9OzA2OrVHhCSdWiuSuZ+LL2rdqZaSG5qgHTTpFJBRGTmyI3K+TxHGBG99ovaJyXjhQ7Bwpq
GuFqNPVqHxIOlKGoTUphgvUt99CpwrrtJ3N9IAIs7rsyv4D3EUTL7hQicmoWHWaHzIVfRct/oRTl
AOSOLqKCaj6RdeiOwLZ10RuZGOezEkXBSMh8rCNTKn42fd0dOYops+LPV9ixEGc8xv4mdnjYQ4bh
auMhcIm5FoFe+A8rWvbdvO5x64BqpBRKOLsbB7LklxnA6G7RDjRycaYaZ4zpYfMC5x3kjAsYffeY
b6tXMU0tFtP9nH6GQtjM87wxEzissDNxDUUg2edyF+xscXlNjaeHI7CNJB1ez+LnthKUkE9js2wo
WDBIhj5JFGl+G63W6Vh3X8IrQ6G85bohIfQPUR/r5S3rEId8OqpEdH2KDHkPLEH48QvT+dKfkuZ8
f462CpdCBRjQw44cDyUTUD/eN0xt0m6r5iSlB+pifNjaRva5zEVDrmITNsmVo1QCvVIUwBW91ZbQ
nHdGT4AZSgvtFd7fDRq10JugVRVYfSfCQrW9RuZHOKcdnt/frAVxESjRitic9AzyFDasjognUBtv
TxsQb4n9vMKijLwDZmpujXCoxj0VZqtvpt6flhOo0CaiHIowP+RzNUtRbBYsvTCvOvqhUVhBaPYL
3sWjZJmBN1a+oHqyeC6oXTxjjYzj1qisHfLQ+fs9xz7LYTqi+a5wIMum1mXNnE8gniZIsoVwByl2
oFISKIP5rklJxQZtsysGJx8K8UGdINzXqR/TkZHJVzOMPXrV3cLVbeoyvzSKQdvSSPRJBEuQ2wcg
N/yrWErdNK5OhAWWsAVvtAn1Z4JTOLMtDOaJbXmGIoWKZWDoViLqd6HV4tD/ogwAjUGn3UURQcaN
Ok0z7mMkIOFECNC+W4OikOOUY8yOz1FCowpaehoTNJlZkUMiEt0vLVwS4LZMJrO7EdHhUn275xWn
QFhF3gS2JmyUjE1E5TUmx5zOyO3hoE3IkKwEQuND/ouZIV9D5stTBR6UOG4jAPAs3hU/AlNZtmcs
cohZKCguk4zGHx2F4rAUu5oWB2nj/5VtqxE7d9XiYzh//7ZTLQtI9lPjeEaENpwFbM8BLjsFpsJq
wC8dVky6dkGxjpZfz3Kn4uSEJdcR15FZ9r1sC1Op17u4v2MZzVISmq3DujgNPVRp/BJNTuAZRAHP
h450Si89UYaBU8BU40kwQQy4LAyBzsFlg4aelmQTwNQ3GSLhT0dZGEu0nfnnUFyXviOcK4Xib8Un
Gq1SDAOsCN3o526pW9TXxawtjOQhGiHCRqBTZ/jtzPvML24WE8A0LyWuEr1J3oM36cIXKzP95wiN
4WLAoqluDZT3EWXu46i8DqPoxTPRvLtdE80SNtnOT4bincuOr6B7/ScI5rHCuv6E+z+arvO97b/Y
2RK4MR+LJ5CG8/SyO7ZQd+SeDPKTo+eXOpn7lPAzZn5VOGZLog0pf7uOJDXAC+hp5zxcEXfZ392+
vPg/HdG386SSpvxZR20nvpL103Z0yqCfbgOXSXcZG8czFtO5ake51vtFQUUgtuJs2Mm13E+fFsKj
jFTgDrNDdv9/ndKRRM0cJLU5i0SvvdyAidaZa0bHQF4PQ/WnyonEiJOqNPfvzKXCh1VIxtxWKkPK
8KytDkONG3V8SH5K5afx61BLaiN3k8hIT20TV4cdTaYig2dR7YvPNP7SGVxP8Gqo2YHtEHQzSrF8
sezAgPvn78y80WnMdumlUez7NsR1xO0l9JSxXgem+Mf8uMM9iXZTu64LDG7JVO/y5r7HH8nfQT27
/LR4pKcIsF8FcwFT/Egq1J4qCjv6G/HaXpAIaNWhaMcNJPa/6HRYXvgGb3YMwPmb+K/7+80I8O2f
5aB4tdhsx4RNVTwjrLEwNrs7aYjgTJXmXFeodCs7sLKai0224Pew5payTpXYI0j+cRtinvmNiOka
jFpmpHXA94DnrkcrHb5AZHodcsOs7iPiVsVSEizuIptnfyupnVlCFkdDiY5/Kz8nOB1/SrAkGDmy
KZkIj2zZuvZ+M8uwe8nIaKHZBqQJDGiwFDsgemH5hvTwGcX5l6aijRaVS3wuWAl/+HtJLARZ3wPz
u7YORcMBtrpR7ooeHCZnCDWoSo9TGfwqW+7k7QZKkJJzaJAam2Eg0z+OgHIbm7Pxtt/EqzOFEQ/h
83thS8hXv4gFRdskgW25nw7lFsACMVD6MZKdshA0ia7geu5rqq8RKb6/862lLwiupPpuT1y68XAB
1+m+psjqzYfuQyybCk4Y8sSqGGUf4uxGytxeU1tuasbA4Ie8ETkZILX2619klK1JZRYslPOCsbq7
JG2LZyXw5SgYCShRq2sMpowWJMGCjGpNen643iog/YTOeFhhQeJh8klGqFLo+ctVE6COxQie8nzy
PBA6tsZS91YK4UX8Uw7jud787ikjQaf8oyjZ7k7Pt7hQeAaL+o9JnWfXL8VLuoP9OAHVd6lls9oi
2kbxugCRuclfI1KnlpJ3nJXahwXhmOub8yuq+7UPkYvMv/omvQzt4ztFtOf9d0qu/YhVd3IBkX06
aAUE4b13iimk51NaXgWqEDh20CqJDGphdaZqEUvEa54ih2Kcfu4JZloMgY+AA3wPGKTOloZznuof
41k+5653pZutgJj+o5YvWkqdWkafsCiDrLVd22BTySV5eTpGv64QDw4Lp6C5FXbYfqsPgbJOHPPS
x9lhWPZFKoSHPsCSV5wvhp0Gv3clAemXLBUgIqB+U37e3DebZUbniZKA98CcNW2J1QfV7VXx7vXm
y7kl3dLiWc264v1DooV57tpsPhiPY9pKxLkt0UnSbUk/5fHz85lvn5YHeXUr+2Jo2ROydWPwtFTx
iyJnLWlCDXCXWCZrv/gjXnqP1tC66npW8lyrup9vn7LibLWnugEPh2/Kg0ppRf8VZSYyKATPwl3w
gUP5ETLcjQyfZ0V83UBKw82A8XEj/JqU1uLS3H1hvrZC9Fws7pEscB2r0XSi1Sl3a5dYSmKwK4/j
f9OdrVihkPWS4py4ClJ4SQTAVcV+QbIyxgeCbYnB2DEfNvztNAq+tKtLTvKuOSY6FG2zv4NX8K5k
AX4DVGYlg6JF3BPp1DHAHURst7IhfU9G9ERcgVVNc67mxlIwZpinwUev4qPQpN/Mnb2pFhAEtcAK
DEqqU1wT3xu5yoiZkN1i6veAQ7RMd2htyOIZoWynEx58eUpLxtlqW1VzdVVhVQ3p7P47RPKpJXnW
sHx+OgPcBZvDWNrjCKFgPCgmJk4qvPznHTLq/9XeHE5sFgILwVd7Ychx/Zcfox7MXJWMel1wwKrF
1nGbYii7J0MOzrA5Wp1ZA5fZtAOurCNk1sZvpDdtk9FQdwfXP5DIK2Tlgd1Zkp6u9z8CtbhoFaj+
/B27zwCDTzE8qnskG9f/BRMT0b850SyAhNdpHGnD5ZATQuJMO0PKdk74bZnH1kc8OuCDUOSF/OQS
8LcdHPb8In1GzFs42pIzsppBFdeAgW+WhOA6uFw71aquxAiYMdiq/tfAk/yJ672DTFjCsIEKIYzv
rWuDpMIFVGfVL2dyjPBKEM4eJrHOm/aDmLG9SiNn2JLQrjUrMlitffiVyMxJbyDXME+BvAgz+QWo
MbiXWR5QMEzn32yVwpJtQKuAPbViNeFx8JVXJVDEdyD7htTypn3TMDTV1NMfXfdgaw4GsUf23x65
Dt1HCvT0lKFe92xtMfspF0h9DnW5dkZ1IauXcBNSMlbbXMWNf63DbL5dfZeA419EPpJwBY5QJ6RD
QF/+S8eR1xDDhuEsBS3D4BekRM0NfqBmJqBDKIg0mC1LsbsnQUZX+8xZZwUrIoRbVOV+etE6APBa
fj28ROJ+c8NBf3wOR4xQZMlWYEKBe7wp+AJHp27tnAeMUuoMBx6uIfV/Db0kVgchBXZL/eOT2dCb
LVuuPLh+i2rQFUxC8w+M9GWpNiS4tsMT8N0rJ0OZx3S5V+kdz+iI+R/NnB6KfUOvhjRuy9F1Gm3U
d6OcZ7c/TY0FpJyypgIaYjVGXAp7PxLmnDUSxcdYpcXdePwq7qf2k7XUnEd8uoUugogq607DnWPo
oMf1Yv2wtqRaPX8hVIMtkZraTZfKM137f7OOi5H6SP2kwpFayRJZrYOwuRs5kUl4+3nRqtYbaWMJ
nzOKdo/Th5Y1dhBN/BdZAsZ9T8+OE2z0kSsftpoGiMHW6xCWLqaCbmrtP4Oh8m0G5HMPj/S9Gpq3
IbqVmbcRTbWXckXAAYJTdZrVRhrQhl8wy2tht794iFIWES3RTwAj72+D3fg+esF7i9+oAxB3DtAv
FV813jhx+lsZt/ZBczdUWajMynlmLzY467qwJIwbNZjBZrfqZlSgD+Uw0eb9EKtLnBf+Fv/mb71i
CpQCVxXpT7qtNQm4y43/yBnRsNVGPtilT6hbVn4sKItckkE2AIL2TISSrBAGWTd/yrad+gvCY2/1
CdApRQOVAxNiiKh7ko5lPqsLX81A5FyMnuKl7czA/M2edkgVglsbkqIU9ZSZHQ3bjXszsl37t/2+
bkZvK5BayyjkRV4ndmU6e5Eynp43BcYKO1IP+TMkhSJIlGktNkXWfyeauwbDF1Y2o127qcokYHd5
01JFv108amuPywyyLcp3BOHN2oqPOEZtTlxdU22PsMQqUIiB/A7SGZCoogpqySttFxx51JecFMZx
3TsNlatY6hIqbi0oyf81QDnmUhyqko2yFhrnjNvhgIL5OPOzCs5awNfiPJ196dqAKF8JrF9gZ04k
h65MBm2pE7s85xLLDCezI7UgthNtqybzGP+h3DQuVWpWYm1T4Mo8raOCcn3aVPmQyaaXqLd3fTj8
fEmU/aiN7zHcxRjYdwU/Ih78LDEe2TYnPTyu3wpGxVhlXnxV4Y2khAOWpEEYAokrwsLvBK1Vs2Dj
1qMTTJ+h/rdk3xvvmFMwtMefOJLOnoaVwNVRHJHBiaJUJdw5JFWVTfjC7NNZh8cnx/NlzjEMTiSx
kcl+ceasxMx6NEn4WE1iNMZWvJOd5HiEopcCyJ5qQuHxDn5wbi26vG+RWNsRzOVjVYzPK0AMZKNB
SK4YZ2RaY2TBostyY1bS5nv70fk7L3yuTBM1m1XmlXidKAyGCjt5zkct3A2IE0dyn3nU1unzHTPX
0hEmymuwDnEVomCxzXwJ+K2u+3aYzggUA3RkTNzNfv/JXJdCm7FjGeiY7Gol93FrBE+KrCLxjbA5
M0KSSvrr5qRlGV46FiekZM7TMIM+jYq7UNtSOtR/GMG8XnYP3IvnDGlPqGDfGF126z+2vhqVg6wq
m0BETjNmMgSSlSv9a63aEQbTSMItnNkuqnlyuoqk6YywPvLEaFRHZzgQW1NiLH2m8+FuFqGz2LMv
gNjqN7wBfCEEQLJzZn6b0d/AYN/llkiJuZ98fvembu5eY2d+s1CB/7Y0b8MSaGMw7KzBHRSYQiNZ
Xx14FhrdnoJ/j9n5zg7PemaQTeKkmLRsU1B9lBOhYyMg+kvrj3Pc0dxWiCVUKdQ+yt0a97jfyfzm
wlUV58nR5HHnzG7U6Nka22EJ5IhjFTUcrZAPs3EJIARYYjzwzb5xvN+LJutFGOrmqxtVkQkHCWhb
Y3UFag8YlGWDMj19MLPk+3WWaIRUyyhbacZ4LDIAgudyg1zI41+t7AfFDJMNnkyzMfCb6M/hKs5O
UZSP0nQZQY/r7wUCy9BmjkdI9I9hvXeyIk71PRN11dQ2AgfndZvPtwT8/BxWawb4e4HPu6U6q1ZA
/2SrK6BP3bKNfHmITfWBEWlBtufcfxd/dmIZkDvNag/4J8j7yYcQTbqH3mvWfKbyW4yJah77C4KY
AQuIWejL9kxWS5N6tmHnO6HNimwFPtXt/7UzWSub6QoSb8MkJZeNF+nkAB3grzjLzEdgCJR1zmCL
7ygXJ8PnJYM4CPCXRkUfdE2k+4BNMcHG7oX02ryWV4T0HNFWVkbp0HMCOg4OMEg4uPiBcPcieOP2
CVPSM30HzkTm7hMlMamHevoSS941hsG63/6fEcbVujAyftKM/MGMpXtivc60g1sBJCaAoBYWVehA
07j/OaQ0zsQc2l8bN/5PPlc1o7JbRkgRnbMeYVWK+0aDx6HY3zS0FWV2YB7rW/SjMQ5O9Y2wvXQE
ITVNEeRM05D85trLR5PKiouiu5TLDIt14d4b6N2MVoQkqVIO7tpc8aEceToyWJz+AU17zsdq7AZy
8DIHf8L6WUOxgnPGyocCiQ+FTB5ym1eTgPtKNcmZN3OCnkQImUMOgAtww9YghxYyWuZ4d6FdXjcq
pEsmhiB24JOCx+UFmG1Iob5ORQoydP54SvnArmWDPOJwDLUrDFgzLYgxyxWw2/leuNMZNZ2F5bEX
fldPXHYrqUVeQAZt4J/AFyaInDKWMt36wBvYtu0jizHmK73t5eTsv/OWtcI0Jzvm7rvaYDEIoO3N
aNfiRN8e0YqG1nMdZCnthCQ4v6cTyPgHdADMVhVA1J3TXUx89uPIID/CxKARfQSCKGPgohUqRCRK
Ogh6z+AWBEU9uJtcGuEJ9T2Ros/57aNafDS5Uxe6kaujqE9p4h79GO03dVZtGLD1yS7zT43K13wO
tPiVRxRXTQ7vLi8UYPwVBLK3gWRxHrTkuBW6pb4AFm+YNCmbeb4Sb70DLW/h8bjqRfdU83bGEj7L
k5EqneGUrsU9TuAX5kJki+1U8b75e0G+iDMA1QtfDGl1u2iNgEwltrQZ8JJyrH+8knHI6l4eP9X8
tPtHhvT2U8ZiAeCQuoKNeZ5vrOSRArcYfT3ZZFvZpPcth2SEi7heKDwGtStcWwgW2CvltPe5tRoV
ttjLMGcq7v+RQyBkCyqCA9S0rhFQGhquICv954Y7DGaq/xz7Pnc9Fvz2V3oh4X1RbybCC5rKoGw2
d8ufGSG45aAYmUC43wfoYMamOmWMbMyQsmZmEikbYgEdd9RY03ZQZWMXRF5XIzLJjuQcgm6wlepN
+y6Xc1hZJZBO8SQmeJePtTJQJ4Pa8DuXx8MtNeH2MSK4wYigkRHEM/ujeWK76W8ZA+Xb1Zvy2264
md2PCBhkVdpT+HiJBd2MAxJMdHUzjAbulq9a0BKAK7awL3+aEFWPh/REiI7dA82jf8A9x2T9lgq1
DovbfMKvPDejFZrrlI3bN6PTWHqzMD7KXk3KlPn5aNWE6i7lDzx7jpWEItQwowPWC5U8JKdQAbDd
Li+E1YwUGtO+aXrk052e4VPmu+vVo+639sRWengOD27CLI3wYp4EGyKKHffW9/rELrgG/3R9tXRs
Fam2RkXPc0+284FhMg40tY8ZVExF10gNCv3zzw5jnZtKtwnc3uGbYYT7tIyI87QuqgDSn1T/dX2b
jaBPKwUn+t2mp1a++xghuZigIUshrKHoW0FCWeuuyemcFJvmxb+IHYl52nOOm+7Gec1bsOAU537+
jzn26D/eK79cAYZSZcon0WRrKju/C8uotpCJeiZtDexZqWEjUyp1ysbc/JhlcjdPapiGKfcTL/Lp
HxVDDKcB25CGlOC3q5qeHC8upegoNRWs+pWC2wA2KA3vrqyQQkAK/nielXLPePJKukY1lgmSq20I
ZUE98NMMCBVc4vlnZ73rVQOC7BfqQRNtSf19nPRY9IzPTyxBXAOYgkpeYp3bQbC1u6UGpkKwKCfu
eMz2Tcg1hCp7N/iix3uK2wRlHeSyv5FTPVJnnr4Tmp6t7i2fAn2EFitEhp1yX0P7Nv4dn8N2XUTE
vzoXVNrroZo8QO2d8Gz0GgWD83h2/6MFzMgcvDk/PfQXKD7rAzxScfLcHs4uYra1Yzo15eSut6R+
z+tXJQ2HAMhVGJj34aEGavI8hYgbkdS4F0xawjMOVTVVpno07gjBAbtLMVt8bDLVl1bU3FxvsJjb
LwC2KGipiefXYHOWgrYL/BK/5mh6nhdxWH5mMfiu0+r7XdvFt7Xnogngj4kyyntuS4mlPsG/lRye
Y9Qdo4pn11c4UutGPgs3pqa7rar4KYe9D2Sxfma+8YXr4qW2LQgXPpXaSqqz7JZ25XG8lMKeggCL
XeX76ip/ZIh2Gbe3qYu1I+qp6/7k3kN66Ilu3rO5OpFag+zvBUyvXf+yAKc4EsYuv3ZyXHBvqpS4
WC1hGwmtPrqxSEjsP7BeZoHlJZeO6/EPLZumr67g11BP5dS3v9QYxyhXO/IunuU2D/zHlZ3GPcgG
yDVLbTDARdPsLLuQawrI5cyD0RtxZrxXmEjm1AVo6KGONGFukZHdaVRg6+Eor0hHEZrsA16p4luX
8Anix00JPO2H/dLp1pVWiYWnMNjdjDnZN+uAV+ejmt/5FzzTOe9CUNzJfKqzX6MTwEBFg2DdXfev
KTjhjbxHEgGmfcGsKHGbVcUBMrm6hTr+McA0sB3R/tcxmtFRK5X7Si29uXS3pCyTUNd1jsyA3Cu3
jITmOYiD12gkR+cdaOt2LEBKpplYd66BIvV2185UuioJJydASWl8wAGpWgCZzAkduhgdzoMwAgHP
raHpG1+q02+/opdMecPw8/axxgEi9W6mypjVdPZ2AraoVw8svbU1tMm9lteXHcih1MpEOwh6ghHA
L9bb2ZdcEmTdsg2phGCIz2TtTOQb/qwIVAGqkYThOpf//1ZZgBljZaL3hBgVMo/xA0fiSy2LFecm
5igMZXXbQSunYqC4GCD5lct7zvo4UlNHDR7apJgdWc6oO2PNteEO7ajuqKWzVFO2i3P46Hy6IYWw
s16c/5VMB3Avm1sSfnun2AKJvaNZi98okY7W2/k55cyUT4zdiIb2SoUHjyQMJx/mmcy363ko7Po3
x7Wi7sMLhnDdPcB0g6P+sNRdV/+3+qhpg5OBfher3s58LAEfnYxEZoqgvaPE1GBx9YQ/KroOfFkO
x/bAa8hsaq4LwW1WX4QhlEU9TI7rF+HuPWbKr8uCcLKwGKPGD9htEUjbI6hSIk0n7ba7P/cPnYSv
JmJlQhL3lk/ZDlQpbN+18R6rSrXodlRs5o1TtU32sX7TbQ0xOhH2Bav57HUlcUwK3rsHwZBpOcL4
ptgRk4zIP0YTQ2VX026bqpK0ZYxBDoe6dW9h+yhWdYEfhrtJ6OzVq9nWwz4SPfgpG5MNiYqn++ua
3viPWhGeMPnENZwOreEiLl6juu9EjtCXBtbObBAYMg2y9gXHar7+1HUTVCniO+Etg47GbCiFPjyl
2befupVapectBzIO8iXPO1E+AzN0y0p8/CqK7bNwRl/sPQDDIy4G0z7YWpDfq9M2ru4lmjO33Lnj
+qvPgOVIyLG9P3euXo5jXWqg3NYN9NDAYU0t66VwEvC+zc0qZt0xqq8bfHfCDw7ql/YMU9LQdxAS
4Utv9lHWP+6bq6vnAR2RiW0OOzbDIr75JBzUeZuiUoD7nrKS+TmTRv2iCyS7l8x1mxLtjDIPFYKt
1WXI6KHnqCIDWuKQAhue88fhQwCATfbfd+GyMJtTpIaFcwxqszUn+CrqP320fknJdPh0+OGuf5er
xM08ff0riG6HEjyjR+sUYCjRubUF0ske2qgglviB58JTz4U10or20oov4FpT+C7FSO22xdb7nC0b
/kF94usmHEsxIrJGDh6q20NHjGFPCC6w32ZJKftbqZAPb9aFRbktNwduPUyqRju5412D31DXkERr
mjS0TqZX80fBErSZKtDeSPKlGcgGU7YP8s3xc7TJiLZeD9ahx6EamR3xEAu/jf+I0mjCz308r5rN
21ZUf5EYKYFJDki5+XrqUnYelaRL+y4+xLyA4WykiDvf7szBqIvC5rxKg8idlpq/JoUhGUk/vDK+
yZh/qAy5P1nSWFtGcoXINx3PyT5u3d3eu6kc29IJl0Z8hbnrKYTwSPy84/e7GTAOW0kPQxa9n0Ih
BX9XSFXKCVJsdYyzkqT0EhudU3wif5oqKtzdCnM57NBY/kJ/3aF6sn+S3KKcbN+T/NWWA8yJna3M
GubDld7+3NsLEt93KxTmpPwtUGC6FqBKs1F4KwLBJk8OdyZ/sAofpAODiVU3ggms06mxibolkwT+
c2Rd7L3jEOzzsxlGCSq0go1ck55cuB9Hyqd5kQL0UTQolZ2r+/1hM1n55M8ehtY+GhGYkV08hVJD
ObZZ54QpVA3YN0ul71hdhjfnmybeyYk8uEpE1rcZLTRBfUE6WneizAnQXAc+sm+37+TNnsHWGPBq
NNHB3ppBP4O8T6GqNn2QyhrCqje3+osf2BKagMxcUfD9G7r7CH5gO84Hin4yNeDT2rPviS4Hyb7z
RkdapXJvdYSxbLLosDBsuxTGtNop5H/dCOtFGZZ98lffVdX0HXRgqNgd9C6E7M1sAGyESeRCon53
N/7nIdlxtB/MQP1o1pdjNeckSFxNWVWgeq/REK/g0OvWij59CXuUSj823VO9G7q6lLlJVzY0b4xY
/vE7TbxEjQXpUJg7FBVLaZw0eBT1Hnj5TCHeCD3AcGKC7hrukJVyoZqqLh2o6CorrcwZDLji52Rw
WyQJRUwXYUe1E9h2R5U1XRsJXzD6Fyh9zJmWHifoxbJH+p8Wz2AF3ZouHHCmol3f6/5Qzfvkn758
eer7zy9AdEt9U7IbFmRJk759Vo6Czti1lUVx4pjgXqZ9okj5G09/WD45HNs6XB6E2OJGBHLBLoGU
96eKRjS9d7qb59jY8NJcLTxzkxZW/vXRV6ijjvYWXqBKycmaxpIfdKIyS4+Ud42tPIj17Qbf6Iu2
EI8SdI44g1V+Pf9I5cso9qfqzpEcWT6QsvFe7iorlBDzZQAzI31WBy+k8hvoIJIwGWCPlUxWlxxH
Fdogdjxvi1As7Pngr11Wud0N4fkm7AAG2/JYcumxtXc2tokePCPLDMpwEeJRxHMqqOwWaI0VBVam
8QMBepipBRw7wLQgHiZ/iQyEI16CcqlzaTeCqEJSzO9In6XZXLAxZHd88ymb4Ix5Id4jD6JatDhe
HYvAIwh9IjDKIyWH1xag/WnOIR+9gSsVRCLnxiDtIHuqAk4S9YmBHDAb1jkJ2UY7F1J7625vbQ01
Z9tWw6wmpVibzA8II3eipGtsvSq2YQfF+aUhTB3Gd+Xbj75KMIZ/0mTExTBuM1G1zMdnkeyw3WFi
yMpDWrVN33vTtewGdQNbumZ3p7wLoBNa24zvOL1H5888DCXFccWTNoYO9s6KyUvQwr+kCrHfN2ZD
sq813SpbURLORmaFdLaktC8fPY8Usqhx0xmxEhbbYieOeFrXWHt2l1W58fGtVb1NgZSeXBiqqiGG
eyWZiLZLImjdQ32uAX3op0/lJgar3txNMDUwa/3szmLyvYu4gX/k1R8lNkzagco0h0s+AhtRP8I8
dt5iCbEsh9ZaUAAsGHzmrMdMXjcjn9hOAFUxUzcGCkyzDf1egOtJMO/kH8U87JDM+jtCe3pvGJy8
Gm2Q196oOeRwiM/CurPeleAIg1f2RUXEamUUYCkwuTUaMxvsGZKV9bMad+ZYtLLc0hwLTGzOatFn
oEjwuXiOksSw7dbLK7n0oOyOOJKa38Zt1pYwyo7cXF4kPT8z5IjzF1vAO8AUBFJq0NK1C//Z2rZl
+XYBX/vhCt08rbaGvifj94M5+SlRF/03hm7XGcSIXw1pZe051fKDZpgnC2kceu2OnEQ7bslQBRiv
+CbAfKjY4+vundUpGO0OVMV3IaBxwtc3Uu6WTCJJIRhT12KvQpUnfl7bu/PQZWhOOjzfHGGLQcoi
OpqXkdyuk5UtJv8x/lGeMkY7VTJw/sK3XFbrbXqd3+cPZ686F6iSbrnGvA1xVGe7cyc7XA/jFjG1
XoMYqN8hg9wrEg+eGxRPx9HtyIizX14WJBIW6N7xLPN0AIDR5AMvbbO5mGHOPrikg7yXhq7o5VX9
tUlJCrQVOJ5eXErOlLswt6iodOhl2kGSCOLhxZrxgv+s6+ipP0B1kZvEBz31P67pOTRfmRCx+Wyn
uLaaPlX4hvX8BdFKc88NzdxvBlDgfW7F/OIpanFS1O0A0yZzlA9hlmqxvCGtUyzdLhIrryjDUnH4
IA62bVF8B9CqXaOT+ybpyPqF7TZjwBTE+Wmhcs7cImUtG5OfXuRaiv5PG9WVLexp6g+gsfQheaZT
0Z8qsMsLIvwp457vrkewGcDl+0npxiy8JHqirS9wO/o0UD5iQlFF7YtOF7f1OWMvbxOuBP9Kq/Lc
QfD6wuoJLQd0j5oJMfyEUx1tGoC852fWR0PruDbuQBlqfmsLGSY22zyoyabeXsWPL+E+hyRB5uBq
WbOe2cvlHXYHEaTjr4ma668ZNb2RGD/j5x7TPx7p+t4HQ9TNHsX7XXaiSvLY0jCq8DMIY471JmI9
BlJGAlhuIkKDVSzY9UngisthBlRCTsJgZeFmuuQBdYafSL17UbGIDT6uJ0sXCZ/4aYnrPIGPe1iL
et5EH7PMXWElfJN7F+oj6uGe9QU6eb5a8NQwJ7CbC/gNVqmXdxp8nQtUf20tep8BN949D3ieTdar
4cSOZ0JD1gFKSdPkI4U5Fz3WnQ/jW2DcrOPrlHlYCyiD6/GQ7LT9hXRXJTlLV9wTSlVr2DxkC9sQ
oyfUqAgnKP1L6NqNsmAB8lrvVdrUYGp7HL6mGdf/G77tVFBW6rVQwJ/elnWE+axm8a3dQ+5Brgat
3E22gq2LSDQyjRAhs/7Pi+LFgwfY8dBK7lEEuj1SeMv5WBgd5y39/05j3C5kNrw1bOrXd3ZhnWAy
0bD2A7U0DgXb5zdLiVmqZlng6S1zDepd0aDDpYHGQxaPppimDSbu3AQaIvc7XL6G9f8dIrG23cQ/
t4t+uXAAcZoewAebQ0ldFyspwUtWNQlTJe5E7lcdzfyZxoINL8gmxtSt43jWeFz7NJTHwS+N72Zk
5cX4DZCUW7xrkzUSvdzttcdYU3TPhVKtZMAuAEc0D4z5CdGiu+TB40TbApPl/6tcnH3TK8c4ryH4
ECuodLHGq7bLN8Coef17xnFGFCe0dUO7CZk/IYvedvYKlJQ2lgXQRKYjDPg5fTsUbxcOxvy5iD2Y
Bt4tgGwJZrILk5gUR6NRdLYhpuLA/ALrYa4RoCUSHRGi4RDU9XeAH3g+S+eKdXnr6Repg9W1RdR2
p5CRezhdFf39JezUTtm6NR9BQC8dGUw92AXxw6i5JAWeMvNT06CLAXAajvKicKN/bwqy5hpyaZ8v
GAYAPVHnfcDGC2I6MS1GF+NUeSzFe2ycoU+qLXekQ/KR31S6TxqrZhzGHg+eEFgsgihCoFzP/1Zx
bQASiym+5oVanmivCiEm5jDfS/5bQRa05l+T90U9s1FTlceYtkJvCYAkhcqMUsR4IXN2vaQeyWrC
G5t1NTK8oATyjNOQ3xpTGPcu5V0/EQB9gQtcR9WvBTiANz3vPqOPoov7HTWAR8yVVac5vDKZzf3P
arAdw6vvEJ+YzpBgEGrkqDMd4GtDyUg8icXLFmMRGrDmBY3CVylW54uZYzOKwW+U4puhu380yK/y
BjoKFxP5H78I/dGm/cB5yzZtQ3sF14Y4hJTI01rxRYI7D5LloZwqzYbZdo1fvbuVQNVZaH5Zgsyw
6tTA3cG67tUr0/zxMy7EnqT9jF5baZOO2KlS9EQDqOD5hVRfB98feSNOC2lrzkNsc/1tk/8/CSSy
PHxPxzm0at6CuFHqXE6HDSCRF+PaF/Rd/QsVb55oyzyGR6jxrFoki5Zi24rSMVHfzO0e7xt7iN+i
joD3V2ynKCydOMVoNRjoNkTmDrzfjQJusaa17B1jz8apqQZlOKmgRO+jC18yAQf+qmz3eYmlJq81
95mXY2irH3RHoLQ27QMNIzMFUtZVE/nRVkY4LTL7sXv5LdxnCxWpMtr9In+C1uBNnJ3DsBKV3d1N
ztfthfxHVpx/V7t6a7Tm9NphnHrYn0cB555GeiXLGkZds7GGrgMeVuohwPuqBq6y16d3KvRnFKfq
ETcGJmgP4DK+HeQ2HpPo9GOLgR8vhqz9KBfHEnUJXUbEsvqLnP/Y4+XknZhCcdMgwH+V1ulbkyrl
LSgYUtGDhOQMaCdx0vrhmkL+Eb66yc8pxmjZuAGSfT9GUAmNoJunZ5IwecjbsvFGPCWDXhS4f3WT
QawqV6DW+QotOr9BzppLDV/XdJtfkl9eXXJac+saJvPGl7OZKM/sU4C2uPwglIZa+mDW1kZkTKYQ
+GXXr9BazTHe2w2OrUSN8nxmRYKUj/QszOoDr0f3XAeOfDZJNQs1UUke7s2zyGYEnHsPwv5dHvba
OzQbrRJpE8iojLlJIpYGNOkMV5URAzLZ7PJLvh6lv9vD+pBIEZgPq1Ivf+4h8ofp/663izcEuQWR
dqij488dmsE8xxZz1Q+QlBKF+BOePZQVM7hCdZgTUnNzwz5va86d+5C+3rbqwtLrxqHnAZwWJhdC
5rFzgqkSHqOm+Wc0ytK2HKR1UObsh4m6PF0Q1bEoMIcO/DqUkBNvilI9g0uc5sBSNGmhN8UCzqKe
rGAZzKNm+L8pn5y0MVSjEdK+dsIPaNVho+9MfO4WA5TAs2Rn+WU/PeOZFNGEgaGdOapreLL7dI+x
EpujVvW/8ud/X1h8RlhObTCENy20svLhb64e3Am/53TTS1jByj4fq+j0pWtg5vh6tnUth30c2Qju
lU+e8hx9DF2B/jIcEom5pfayTbYVwuWAE+X3Qn8BQ/ttT1fiKTunPOO5i+k/HMvnpfifdOO3ku9B
Bi9x0hc8qXUSc7tl47GE7munw8KJwgz1GJZvt1WQv18iFJA/IXavfRMAadLXfmA1NUAJwGBg0gtl
ksVOLzI7KIFnrxtbXfuRa95lSfyvGPoMNmVbtQdehbaLgIx9mYOFsrdy6UUPn4zZ3n3GopbE4vVY
hFOtbMmjU7tP5I1d6SsgJYgUKa4uUs3uyVomewOz90TN5WDa+823WTSEeAceG3pD0ldepsLONui1
6u2+WSDUXz+iVjE1Td1aU7shdj6+M/cM4mb87x6LdDes+v7miAOE+H/p2PVMgBR/8bAIpVZN8xMV
RVrXlZlgRp0S3cnWWWbvKs4+cOTfcUPbtgUYuu/7sU6RLL2qF/cwQyfGYNfdI8YJAy5qTJWewMEy
VGG3eXYKg5Z7ogunWQoUwhz56PKoqBj8CQBCYsTEARxtpe1UU2JK8hlbfhaaDK6zfO4EpoGEzRFR
tf7XWiNQ7qPvkz881Vecqem/Skwm7iDwvqP/qcCpjHKnIELCpVfYeICeBnZsd0Qcl0xOdgSXLVlb
+NIKrm4fHF0UZLBV7DeAF+p2P+zmrP6N+IeOtg5oMHEm+7CikY7H7DCYPbAc4lp67PM/7u9jvSeb
vYxsc0prmPbbYkAoquB8+nK2NqqplPF3bzGph9Mln940NxQhQFRwon6nJqBHiX0nXZ1c8xloYikk
QkP2lP5rNbrjBK41mJpz79rk9nwENqZvjPucnjzl58T2EhutpSCv2NSKPd9O77AGmg+z6pGMxER6
TffVhtK27MnLvN9A7Oebzu+WCsdZziGy5h+4kvO+8TOXTZNC3TZOqtL4AfdH1MeyVDKzTbglkC6m
chYmNmL/UEKB7U5Qw7gjxvdxHjTt8ZPaDnALOafPUMhugEjMQG/mh0fd2itDVQa6DnJJvr1+RzoK
v53iFc/lmuRUkFN7NDx44zIhf4Vb+8h2pycX7aBhCkO+LlJ0yY81W7F8yMewUeveJj1xWtx7LEoG
oGE0i0RkiOh8kbHVZRUecBUvkm6nqMv/xGbkf9xvp1C8cafgHETQzKk8ZC2DXQWZR75PCbJ+wGzO
r4zd/UWgPP19bPoymn1vKyE3drC3ryyBbGYA6DNo9VR0xQllwLJ4kQLoZDA0ZBrKj9f1R8kpRhNL
sTLO1+AZ+9MatNu0KuCHi9EAUS6nnlFunPhLiTbDOtgnZid5ix+Cd8Oyxt8Au8+dfq4bdZVTgNOo
uQ99Ok4SOxiWlu/RnDa3RsfFBZwfIhgMgxJ8AzGafn97DKSr9i6Nhj0Jskn7AialO7IjlfkkOBwt
gHiYnTLG7QHWBMqoWx65DsDSSb4XGqKb911llUVmif51499gZq8wLZhAr9q93xkYykgg8ZkLhntf
ysQRGnkwOeKLb/LCgPOwOCvsk9RFotaQF558aNjKhl7xcF70lWieIwTBdKP5uFowXZ/jxjGANgKn
Mzy6YtTmVbGyCeXfYcgwp3hg0FyQ7FNtKclIr1AdVnyP2kExzML6f2+crUNeuRtY8GJfF5Uhl8OT
6QrUBAvgKlJWL++0lFqutQxi55x2gKkQdCDr4VZPRCdTCJ6XQ9nS314FJ625/QKrJVbKsebkub1w
JjfyvfFePNecqHrMtq6UepCeNH1HI1SZS3Hf4gvHoXACOOYwvdpfhKIhyPLtjBkgwCCYQhRC54FX
zG83avH98qqgilQ3h9N966oLEcCr9qAOxUOCLLNsO0AbYArOW7REdrYJdgGF1YpCTS6RqsgjTel2
SdjwE6iEQN9zf+NVmE2cUZ9I3h2VQwIdFmt3E2FGf16O/1BTBHl7jMFFiv4+fa+RFrykZ9T6aS4T
Gk9HIbu6GARvRJ69kZU0CTDERvOaycfxtu9VWAdR2OPf9FICvm/tTz3pdetq31gvXPOeOcrlnuR7
aNNEX+WUMwWT/jo7kqLVwJvxzY8wSQ0CKE4l8TADCjF+IjqxUoGYf1YdRso086vpvGwpiJcIIPRB
8KuJaWmp0PL0t4zuFzvwr+H1Rgi78TIqSMXCVhAax4+0Z9hAF/5A7Iw4r5EEn3N4m7Rk60ucblLJ
iPE2OERfwN166mOYLZzLu9XtxUdOJ44imOYTYkMuH/VXZ7wUVpjWuboH6AkNA7qoNdo3T+/CF+DZ
rv+9i0C32wHf/UdsK+EmZRB+Pi1jXKhiQcwMB+DmOKV0bp7WbmmCn3ranijNZAvPr7O16YobXDLV
jshnAruDP/hF5bSB6r7N/MofExzD8HkjCJzLUB84Ms8ACz5vwGj5Q6YVOsBvtidB9WZqP9pcFbJo
esXXatK91nImQBKTdAEd3hiPQgFl0MdsAWsCcx+nFMFldWptlNYg5idS8YkrYyIc1KSRtzDJKPD9
ZEorMYoP/KudhkGBOY277p/3wTnPwS2GjgXr/LREsT5m9wmbPmMkcCWDz0ZEff/e5Vpf69ITAk43
/OGggJJLZObfyoi1aCLqq5rRaSKQbmE0/vMR8Lf5b05kNAodcEtpMx4QaBMRHueBxwE1GCZ+kQsi
c+1UUilfndKVhp+b5oLlBbPx92rvo5ELnqLxBbVdC12vIty6Tz2o2Wcn7nLZQfch0+avbNV9hPrz
dYWigfHxSxfzR8YdtItdDOpCFsjc+PD+mbdFv3UI8tYBPqf59/07wfILryMMtt9JDyMH7UeHk2Aj
xuyrUE8hCZiKWCNwmhQwDn/b5nrD7S5INVpOQDmM6QiC3WbAj2zfvkMk0Fqjjw/hqS9S9zNv5UhO
Yd+CLkM3n/j/5w0tCpwitiDilm4FnOdKbw1SOmY9lD7Uj7TyLequcLTIeSVPGTCVqR2EKDNJjOYb
KC4ObjzHAtKkjC6a+4cF4WWEyFUKQi4JTqqadvgjUxlO+mgQYvDW58TbfDRZbOhAsLfpD/pwTix5
kJjVMhJqZXD/vfrU+lu+akF92mfxSUart2pVP5pHiY6CiIXQGJJOqncckTKcWOAX0EusAU0OmIkR
IwRbEIh00pBU0gP6B8oi+pL5Ro9MDaUQDFerFwUsTveC0k+okZcRfHt0++aCwaD7iWp8aZHEkZPS
PJ2HqlND7mB3S2/LsZqDg4kevGQwgZO/RK3+KDra6/cIucdukzgPriMvAOE9/FI+W09sCwz17oSr
Jja/e7MLGI7JQgaj5LpIaFVz0Qnl9TM2IMuoi2X30mnwtLb+sn4GDYHLGjLjXXZjcuVUw0Lt5ujZ
PaSI/vzPu1yzUoAflje6Z0Rgwexq8J4TVSXhbpcLmQm9H9EgyRzhNfdzT40kFIJSNyAQRBif9P+Z
bWdPaGrUvUiov0+D55pixUtm8xf+0NbnnqHWjeAtfLCyeaRqbFRYnHCrFrv8NmKXIqQQQ6XOO5yF
WXOANxHGVt7wnPVCuQXnZ+wAStYbnJYAxMoGUm3/3EY0N1PmIxlY7gW2+V7M1Xh1UVjViSh+gtAT
yEBZ7ryQmDNaozk/F3rIgAcRpBmcjs2M7z6FhryifvwcyL/hyJjv1cy7zrHwbQHuZMpkQSuGSLZk
06bLczcRjQNFKFrEQ3ZHEBKEEsyNJAzb8PY18ffPzWcUbLsfylkfDfGCU5TZidRrkfDdnqcjPnnw
/s9GGza9DwHwNaZvfKINJ9Pfme+SVBRMSGesK2/i9VO/AOU49/QRXaQuM3qf3B4uLblQd4idv9z2
r+Q6JJpqg2TMXgz/EBUlQDs69GC9TX7UAHA/cendtEfB0BuOxWVIZd9AIrfFSptkyTCywgGHC9FZ
wadZzutlsw6QTc/dsHMrVyAJtc69dWLjd58quIRlCv2fviYhgo/pByTwZ/acf4ThlwXd92qVWLXf
T52P7On5kr1HAURcrfraasEYGVYUGitSdrP3h2J9t+BmEPMIvJIhN/I++7Xn8JDKwBOjfwT8gjvb
5l7t0B8xB0QyHGNoE6Ilk+lRQVoWdAou5sXnV+JVNq6PyN3SM41sdG+UKuv6LJp9y3DNUTFMF7fN
IAJP8DaZT3FlXngpbQt7rWt/9/HyNIz+ulT1pgeyfNKLrALhU/dTvD6pXr3zydH77YY8tT0oc0ob
ybow3GwCsGdhbF8Lm5EFdcALFAZh0fkm3xiay5HolybXyUcIWwe32YeKpTFQFVf0Gk46FFfme/BJ
bYM6PWfsniuM1I8IAXE/Do3OKxdoca0tQxp3QWzN9YDjYAVoti7cF4bFnfosIExq5KMGj/Ss77RI
WbGYu3U+OKI3QgUPebZMkmE5ZKNKRD3X7zMEA2j8sgvA68ZMfZFWRGkqazIvaBQSvILxrga200LN
oFKkFYFRUgczDZ0SOyGLTfdtv8BLlU//woG2+MNe1erUJIHH9WCsZ1wqrnI/uWA7oYmso5uKoYmZ
pIqJjpiduIEtbtshxKh3Hy6BAln1Kz5HzIAkBkR/Davx9soLo3SGZtIkqM8D1DrG9Op9oEAFlt6C
0bsYUs7zyQ45cYpJ1CgOvmav5Jf+BodbKHJeYPDcXM64dyiKJAWAINxwx8OdfD2IhZBjIGRKLs7B
zmQB42d3OVFyrC0r8VSh3tyOe+atIiS29qfQNpymHWZRDYnIlSLu4d+uc+agGK2sP3drZwSS6ybN
LVa8KoENOpq7Rh9G2+aIoWu1JVFlnWTzfmPtURMyE2SNHio+HXLLmaTjTUY8AxJzuqzbox3gmHrh
d2ntyGcy+Om40HSDMRvrCADcIIxN8k12MtxW9CjNxtQ1IAbwt9a/wjwg50qXvLYyfnx6ArLhDb+Q
ZwBi6CcWIaHbak8stK3f6x3/DKJytfBQqwhJopTEaUqrZrUcquRuVLYxZGu8vfzSQppaO9eEALSh
cApoLtq+bcb4PvB9/CwwwuZYOPe/Z8qYo2AIhMfrajtT+IR20JqhUWlY6+TYtVenNq0iNrB1uxv0
YaakxLrPIaV6yz4dZ4ibZ1regM3G0lCnuSrShTRze8ju974HdiA/we2M+GABGUMfv2oW0aVViKyf
ZFimDvknGES9rzi6ThsNiTWKxKm/BTLBnZiNzN1j3dYLke5Wn3QkWzsN2Py3P14/RLLCqAivT/5p
5AobOLpzckgksPs+oStqfCnLrbYl+ryE0z5zZCeouvDdF1ZSjdak0pSU1iUfdawD2EyC/iCCOQHK
ijpOzr1YbnUT9w0r/yKTya8iW+yoDFuVTBteTQaG2IfZPrZ0MnNxrz5zre4lEltJjrnWRCcSHFjb
R/MkIEyrMW9btAcpaJG9rNFJcXf4/+jScENitC0C0e80HxyubcJ6JggQf8nVeR2YzJRMmsTi1xb1
Vh66+y+EtrsauuZAGI4fuxeDAkRloRuLm9iBet7mJASV9tFwymBei78U9d35HVGHo6xDzqeVR5BG
nLr4Ik/uo5ZqnMqTdeoazXJGwCgboLF7VRKpjNjVkUftrOviz+mM+GFoGl1jp2j4dePmJOXgTBo1
8B1f/ALhPlM8GlHM13IsIjEgJ4yhPCX3CpsLQBsTq3Sv7TrBdPl9i6oHLyfq+ZF7tjL7gtJ5bu9W
hxeTUWJY+ofUXJJn0mpIveRk9qLPzV5VyO6Rg+g4VTgrvYxYixkGEcE0iCNSRlVE5f8lyaI14VVl
jzjnSkvE8iSEY7VupDDQCdwlBDs10kitdA2K/M7pzL+e+WIrCYnUgd5ZKh5qOqeXEB6dASbTzZDy
aS14AHHnR49GErLfq2e+mpt0hMlSviG8oXObUlSb9455ZnA7zL05Gcc7dv3nFaYkn/1AJEsej+TN
ocEF27XBGN/2b95huUTZqfOa5z4L6OABhBdQicOrnyMlUXSdcTxZUfQLNNdNsmOzOpE/fo97zPwy
/Ylr1y/qPS2sHnvT7QmR35L0r8jvykjnzdpfYFp4jI5m/VbFA+gtqswx1ehem98wY0XaX80GIant
961Z0UekUIhufTPnKQ8vgBl/VY7x3laOYKmNElEri9uNV0+sl2/sdHYie1iMCLpLLLYh26NHwHA9
3fiiWI6lJ9x/2RAstPMfZgbmXSH0vqzMNOw4PGpyO1Me35d3cFgfNQgFo3/eESUXt5TWze0oOa1d
LcliCKbtZwe4jcidZhDGJjIfwoaZLbLr3Wxby42vcdrZ+iQPCRxXhtFpe6Jf4BZMrFo1Z1Rk2xi2
y0T1syi3xOZi6tkGn9GqhqmYhqeTfR/OthTmE7VTOxtmKSZg5LMP3P0pQeP4hm0JA8Eprxoea1k6
DTTh6j5GBzcoVFe33RcOkeDMsYtF7OxaY5Vya3WrrFFvChkjDtJyMVoTHKHtbVD57rCLcjhYdx3T
Nheqj4EKm4Ggb7npuUy+6bh/ngTcDzmBZnTNjkkAcYzb1mZHoCGJqRzTjIJKmXCE3PSzH1qMmplT
D9GCzUFGJkxiDLT9aGy2x10PXQBWnuVGWefMI+sWc6HfznTOajS2lo5PeQNOBS0mBbUtHbqu5C5x
SD+Cq5TDAFU3CB/MZUeZGjre5t5mfO9devi3WMvw3BuoVDSpsTVsGmcqP5EPY3Iq5xI0a1d2IpsZ
odisqBx8Jb3qT3drRExVVYzqhheA7eqcWcCZGjKa6bFyqAjBs12AL/jWJr9HGg34rFiGlJGyTEns
dl6mXMCUdwbuf5xdt9p5kZW7LswEakeNYZCREULOQPKf1T2uCCVL0hp/P6nXqFon7d5aZKqlVQ5/
bn/q3RS3W+n/o1Td3VqZsL/EYdZFGT+qP9bDuG3CDwjHflTIbnwsNaB3gyz/a7y2Dxx6I4grPs+d
pn/yLW3HnHDahNIlhhSZb43nhKPBXLu1vl6zaWqULpO9Dm1EgVpYLQtBtE4XdwRhRHRUvPMA7HoL
8tdRsEHuOSi/wtbm4PMBAFNA6AMoFXj6FqyEPPvz8L4C7mlINLYrghOFMP69C7lDv4shwoQoXupr
omz62L2nW3H+90GQ5lHnl/FKhE7qNaf1FnnHCKpPtHEVMybuDmjYyAsWT9EJjhjsFOyOzL4cPGl+
OLtkKiQwu4OB0m12luroUzqViCkL156XvF6lDmtgAN3AeMJCEktB/Prx0w7tGwKTr6IjvQcpBKKz
+Fg1rK+C4epJULvkXm0gUHGyUw9FQFk9Ipz4owKgpdpefv5mXKDAY5GaxE+KKs5YOrYoslE8yh28
TdHlBaOJBFg6Wiig8qEJTEPuBoPnOJKlul2n0tiEhJHreEnH8Euc3g2kPv6vQuEB/iROv5CEondS
6tojMOnB7TYw9OxsYpirADWO10o+9/KOKu3s0+ZcxjEQHe+NuwOP/+2+aWQChyuWecNPqk2muVRw
Ycl5fA55ZNRHz3ychmSmIxJZTGIMF80AFvwULGg+bAGm2iBY2Y+iOJ77sg2KWPkBQ5fmYbvdoNuK
OsWyTuL5SM6H1KzuQ6NA1LL0sYfA+K1YEg0oki5V9Nr01QGNbstxWQlAqQ6WjGVdomSfWJOixNqj
4oTF4XD5TdnpWhOCOYkPJBC40UMr4KCykj28IHn+QCqiEyd8Xs4BKHq6HBV13QRpebLypKYGP+It
KUKUF3WFXdBYmo6UwpUeDFo9ejweDGDMhX//5XK3sAc8QiDjJgKm3MbjkVjOxf1f7/W4iHWYCoPy
ZAOFu8znHRInSz6Y9+VLzQ3Mcs+Q5Yb9TvsHVq2QbiqX4XpAAVODz0zfdpbqzcoD9nBPxMTzVqi6
EO1Ansa7r1hCv72gfMgrQL53r2hdiopTP+sjX1dlkvwwzXQCcAMLSeUqweE5eNPkJ+A09jyyOBXN
Js6lNv0h7fdLfwE+NKjsFp2FfOU5ZKg+HSQfTXGJUPamXy6sMNzk07z+STAvtAYmT6WEVlcb2lha
hjcj0mtZGvf+hBtX0szdQ5kKt8OojkOaUXNfKcFoWpGxBxUkeCDWZDGAKzMkWYl9T2OnFEuAVaJX
djwVs7gxRlWPc03PYEaFkBP9IajxiZhU701/Yn0/Of3oY3r4QehZjazct8Z9+kk/iK4dssU/HADg
K27Xstotkw2zmS70s1TvXQ660stg3/V8MxXhInQDo2r/87MNfIs6ZGJ5bQ6JAk4mUWSxdOIV4jwW
v0MOmp0h/F2ZFi4uNtDmf1R/7i/LXfQpGLnR8xAm7kMCc60y2CqsKtj6NMnC5NHNNZVL8DZGa55/
GWUOrYTmEVN19IzfoWSKGg3HfUyp4gmCwZc1XLf9wzXHJJsPT+aA0ZHBNiOKp5qEjZf9cTZrXL5y
gyQKa8klzLmUPeynOgcdq9quIPvuxVFtWvTs0QVea138woVpu8Bgo1zH0YmW6O+Ya6TtW06sBbNW
B9HzlsJYtNw5Tuy8H1EnqGBah7uFt7iLDieLpb8Gxv8o8S3X2Q3CUdpnnVFzsqtHEW9+XL0MqxzM
Cjm/T+g0y9+xqjlcyfmD+BrAdD4yA1SC8MaGUzn3urdHROdbNZzW8WrzFxoyAOzQ8tD4OhSZc8aX
Dm0AGGDLFwJJN+l3TdB2JdxoWEx6uSTA0gL4zkjQiJSFvB5dCBvBQ9ICXxPT9bnbrpGYY0FHvyhF
L/Er8FrIFFMhyT3dHOwqp5kZBoTf9lKiqDKREfUQkcwAZ9RkuJivI5+cenz2Ig9vjicA/dJciokS
Pn4kq9c42crbAR0s6eHFhQ+c1CtBcyY/KOui4yhy3saV+275k4Yl4N/p9Gwuz295yltcMPMYuG2a
9+4FEskPHMpH/YvSAwx6CzArl6ItDZ6O3eggrMxvojYbRgOspWw5bAkq1UhKpJmMWwG5Dnmbgurb
oaNy27+gtJIpMBwWu5PdK52dEoaO+hn/Z/UNdT2YDyBrbJDsUI+6b17ztd68bkUmL2S+YR9rNZVU
dEiwtaYeAcVuofceycOWOY+39reb759bEKSbok7R06PEQ8GwFqlfXrhpoQbHHIDDyTkP7r+ji4k3
B+fAgd/7vJrPzm1BjU0TieZu/C8UX8byuJla90ZOj+U/rw5JkAM1O5yEr2L4t+L3QYz4B5oGPGDw
atUsKzbLZ6HhZF2WEupcLh0P/eWMkAetpACtS6neGG1Q7Rpdl59D6Xg9528xeAdIISb8yD5I1+xl
Qj/0Os5bjTMLxxEutNuN6VPav/NapiSMG1MOgyvr2HLgLJyszIbF7DtrIvofyw9fpGGNdUg/s6nF
91xfHOxBA1oqb7mpbloYVmHeKchkgoV7sAwOWddyK+5YXXHc65I/a8jEzvsuHXrDBLZzVjbScUox
OhQQTRJiJpE5oMtuz8aB8N6XdGHKxjd0JZPPyiF1f4sKKyl5I5fJo3wKheGS7KHXvM/0h8tUeoP4
h9pjuJ4ECigrYHNtBWbvp3CCywtmCU45l2q1Jym9N0vrSXWAnkUZBRZ1LSAu5MkB0CrDUfgsRsNK
o5DLMfu2/QawIz6ezWdUO0bVtbKRmJRusD8MaRt141JMIufn6Nd9UI0Gaoioc8APwf57h37YZAN4
31ZjhC305MYF437fgvNZoTvP1zy0tlCDdT0DeQy0hYFED2oGl9x9jWape4bo8P9j1eGx3O7OMa5v
f9fhFFm66eli4IUwI7oB/ZVHb8qI+j3EsPPr7h6FO82t4T4ApFOZvVokxHSzW/9RIsiysfK4R6sM
11iVSaHPexTOb2EX9MQYtO2wgDImr+B5OfcB9KXvFUu3/dSf/2AfVhQhW0HJrp+5sQBNOgUDVHDO
kgVBziqm91HnhYbe7FIe+fM/ZgN2oS0VJ/fHK6Log05yU6dvfy3EbDxD2FszkhdH6DpBMI1/iTdv
ycp4u6+yZS9NbXnuU6LFMeA0OKbbkbrQ44BBvPfr5yMWhmgJadcrwi7Oo4lKICcEafQfKPTLrDps
PxVKdqu7E1HrU1cri8cJFPDnISvTyvutPbY4clJiO8XVEl1fIoCsUuLsNT/3juG3iABBoW/RaWnF
Zk9SHsz9MyTbfCu0W45b7Sujp6WTLvP8/GGD7470vMdQix+elO0sIPHY2np60DvKAQaiIdhUTfba
6fpJQ6x8cSBR1i+adk93XMvDB33RsT65NgWTZogmMvpyp58IxXWvPLEDbQqMZh4o5hexKONr8GQZ
t1JwrCiiyGGOPs8fIarFSzUBadLE7cYMNwDCzwn+2rkyPJYOWML8dnqvCubrpRSz2oupDJZkwatH
xthzJKyks4Hl+jyTw28XXV+gKBFMJqafk4CHILgkh5P7OOYI9TtDWyK/exZeiFmk/4lb4657NVDw
2kMHNPa9dgpJody648sC5+oTODArofIdw/RHrfeO7aZTpfVcg5VFWqDw1XF/umkzj6DlKm/3Vqz1
z4+td81IcpEauJx8Ru4UGb6qJIki0FmbLaEzUW5TGUd42FpNIDId35Mzz9oUMK9EF6vR7Tm0/DGr
a6lZqNVTrFeRRsASvM9i3TeixeT4k06PesbwiGIJTFs17nD0nMPevwS86s6qollNQOGv4HwjqUIR
Os/erqo9E+/QxL8moq8ie6rXPZKNgNU5PCV+ZK7l+7UZisDatauJ12i77PoVayZZKBuAAXBSlXX4
IvrzJqVju+XCU/QVBxTHYUeYNriTnDz/abxA5edV3GX7vbF12P0zQDerszePYF86b6AiyYhoBosF
CLPivedt0Y0zeA4bbZ97EotY/ctFhI+XQpz+W2hnHXwEhOsAQ6APgxd6rLCctCQwAGJTUjOYEmEN
hUCP9G6CBPgocmME+FeqB/06+Df7pVZi4AteJwaqM8tkyWhQY8XH0OQW+rvoX2RmBLGvBqYiFH/D
uTgNLTcm3IrCetLUGw27wdxc0fAib7W6psWVw1cdV3E1NtrDUPBabBogvOJS2wbwz1szg0CiXYwt
FDGOtKJFOIGBpOvCCKomiOcepmt/pdcmoP2jFucwbcAPP2c2+5KdKSU8duARMb+NtXCZi1snse2T
Bd17L68TIQ9EXR3CbEOUOpd8lUq6trnwQqtT5Z1F8dYk6I1dLKjQjgOm8roggtFmfwvMIXPDIzKU
dAWK73lC3V2dbsdqtdn3CuuWEtYS4k0OnRYPf/S4W8Lb1JEnqTljj15n4XRWrevYOgiVclyvJuyu
Tlv63SRlEnlrctGFgIoZafhsFxKnMJahALfxy2eFqdwQcoroRze9LzUltcYeJ3+Cuzj7ww58fY/u
VR9ZMeLwJKsuVszpI42hBUwxrXZgggH5KcMMtHNkLdEXqs40zN8cUS+dCjyK9q3MvQ69/GGHy4IC
YXIKzDtAAYduPyaEFXJurpk0Onq+3H6gDXHcBuczLLbCbzDghRNnzUcMiY3ZrMfm3pSh/zjqEZZH
1kMLavr8ltqteFUAviP1bV6aWV5QP5UdtArLC0khACZTad3z6oTm1bQVq9OMPJWCKVGs8M+lxwBr
Wue1+Sqs0ixuPiusPFTf4+zrCbPPDDc0A7P5gUKJWr5lgJmtwAu/Vb6Z+YUaL7Y8/R8zxsZyLuYR
7fq8nVCS6jOeebFofGrfp5DO2/csT0KGdPbHUwroYCidEksylhx49u6qYHuiCUldUZxQkyULVigk
kG+IGhx7oWgFlxudR7YLeIlFQhiaajEG5+3/w3gFOzCWkwTXc8vZZfzA7OtjPMW5KZCl2BW5KzvO
tFBgiuG5cn82K2FfGXN7ZJa1dByqNCTbBT8lWY2b6Kq64uRDhJlS4BhVddqqmpRzB6hEwA2Mx1qa
59j1KSf7xNEqU7RvZV0qg4WIhLURApoqDz9WJki733ohofGZId/imAZmjhTeIgssKxp3+VIde1fx
Y1XIwCMgttprnKFb3IAo+lQWvWh1lvNelO89i4oSOKdRNY4appnV5uDIb94j1o/XW7B8zBd8wzZ6
vx24ejboANNg7Ixjtk6+x8AzruXDDll1wK4tR49HgvZeuiU9ZbUuUN8l4zh8+CeJiyZfe7JYUvCd
/zfMIE/5ErI87dhYK78gquzex5FjBTZ1agqab/1LzAnIQoBxo+YVqEaGLQWZhfkNjkso87rEOzZg
ci4nxFJ1tbnCR4eNZRm92/XBbgXLAYJS97BOhDqOX7ecU+Fx33kWPvRsXiuT6VaJ6Qt4IU1kAuKU
D5Yl1t8CNRhTisFOTOFufxfuT/Ct2l0ryhkSUfufKGm06XOPsuDFGF8CS9wXWfLEBGyBiyGk7kBO
SLCtILdhZWAUsz+mqDCzUiGZXyd3k5wYCFhDugmDjzbWBEy3Dz8V2AkMd2Gzr9bqFLt2oZryXjNq
Z+CzsN0Lf5/o9qCUDljn8RjyEoV1U2Lu9ls4lnvQxZzNkslNOXGKdHy7osvktIc3ZkP+JWT5mbqQ
WeMWLILBg73pTEONTZT/DcaOBSv6ORmL4qoYH2Z2kK0BbIb/Zh6zwl6jZ4J6qK1onNVYQ1//5ojs
wFuoo/pklDvS8JHYmI2O6HCwcxVny7VFiiJww8T95ykKku3DACYO88BbS6Q0qXx39+XeD1AI1Ch4
NXt6okTFjT3GaYpWvtZuGKreC5yzjM4ODDlfSGEpGu+xw9VZXxbpRD0n+AflJ6iKSfzxxc15mL5t
I75f74UAUYSZBvlkERjRhBplqaEB3wBbuqQXWSYxkE8K5llk5rURHrxHyWXt9mIQWQOrrnNRrFXq
W2SE1hSPGMJjvG/gpwb8aCBuCZiP8r5Qxo3e4Su0u28/4CoTBXrgBvyCi/4fpE3GbXL+UqolYmPZ
uWztCuPhqyqwPdCRQFMfiUciq5YKJftIKivhbNs6bnRp3eH1ZCHK8c31mMKV0x1crWfwuZkbQ5aD
I60exNaGuWOwrK2bJikJtu3xOecemuBr3vp4PLGTZSxrdKsbx/0Fyvnp4XnVqxZj4oHgtZ3uYIbE
60KXy6nw2uBLz4v/Vri+38cDGI6Uq78h2obiv6fhV2T64QiahiTJqSsEHPmC/0v8cI6s4kKaaViX
BEubY4Ko1eluc0D7AvR45qcVuL611JAxW9BBguGJbFRY7W3M44dvIXt3PcBiIKvhfKpWR1pWURQY
AaPwK3DlcU56SpDO5VvbJqDO8D7F+fZw+t89tfPWg9e129TLZPeUW2Fu48anM2xp7AP+Qo9sZUMV
dPvrGR8rAZhsk8qeglEd3Z2WO/8hpEd79345OxL8nBbuynCZR4JGqvuHbFVVAV5mvCxNREX8L8WI
YG1dZlGCDNXIlpHvcG0QPNGyA5dbfFf5PrvVbAlz8qd+IW7XDhAw+F07hHT9Q5aUIowAkOpijBjo
nhvHAIbLIOv/VeROEkGOLTJmNMitTLGmr+TzN58gc397tT1YsRswbO1HCxhk84BWffQFcSYq0+Sy
VNnza5IIZR7xE0uQ8hgah+hVxlEnz8EuDGyGTdwsdp2Jp6E/l1IXrY/PrG0R7E1u1tlJ6qZDKTvb
ccOxi1UchCLc++IJqdVdM51HOEu8QAQeDKdU9np7HHvq3lh/0EtQzw2flZ9d1MZ8vLMwwFZpJLu/
JENgcmkkP78F9blEd1SuzywwyW37oLVZdMhBx2qKb+wU55fUKZcR/Xo1BeT9lqxqy2NhiUCdcc+u
guWcOfkEl2Mnkh7XrdZZ2SVCTpqPTYCZh6RpeSCY5C939qppjbRaGwb0FOt6iwAHWfX9+lITbNq4
f/2PJKo/JYId8l3wfv3hEJrptrxfJPYrwfSZcfqVhQkLZ1tCZ/mAD2ixaYKMb8EJ+HwLculvBXjO
rM4QS84G/9cFSjNqmbmLsfs9fHYYYYWFg+/eJPqezWMbVR/SRcUMPezL+6OIeZbg61s5V+DVUVT2
zm+5FWKPCrtewHgaZ9R/XdWciRtrrWThTWteQtKJsXiuv8SlRuSvSKBjn+8+7seeQ7TgrJhKcVuU
eXsRT0mOh4CvEDidtVnxDrDkD+16PHGbEZFIpxGOvB3Ylt+Xeg3nM0SpdwKD35GbCcIRxPXlkxHk
XOc7ZSiwxriRHUTtR4nldOZgzbJ6hxLgdo6mL/JfQruXbwFIU90tFYaC/1PZrDkCG2JqQQ9qNiTO
8FYnrmZIcq7ON8BvNOxqppqgW5sz7c+qU1M6lmcVesLsYPbMbZaAmN0pqFOfuCSelzbHWYD8XL/Z
bX3zCxafWHgn3QuCOJ1wSKCF5SXvQ7WzghDiYfIiLf238WXLt8DRtf67IPN6kK2aTbrLsVgfYXif
t3eir3O1lhWOvgN1WwSq0n6mUgK1pBjWgioFy72rTt5BwWWbmUidTYrdXO5y6gBpvwtLuEbG+ODc
mWsMXv+nE3RQg8LKKWelgiO5dfPT07jaxl5C9rHnguWB9NydoXccGYP9GZ6GovyeT7CJdiV8ekYV
Nqfd/lCRh1sY1m3XhEROu2aXP/NpobkxVJVwmHCH85GBRCvhOWGmrFTd9+p5lkKZfgvHLLifZ9XO
lsM8auhOg0pFhGCoOO6bHt45k1NPm2iG8HHiUpOT2s56aLwoTsDXccXVlQZmGgw80tV1ANiZod3L
yiWDxV1OkNyUR46lXgr8DYrQtb7Krtc1nh3UgEW3hh3GsGElyTawgfTHfJNsuGNLDG6X/WOO5YtX
07aJduFqfq7wABqr+8ABk1TpNdXjI2N9oBA84/0WhQZcedWTJhbpVLEl8XDTNGFuKlCZtEe+D7+D
RJMFEEpVQJD6u2mJv1wvxA46Jgd1LwNjH89jpxoOvrsfBIls+r0eoH8hkIx7RCuG72t/8lsqRk6v
3CJE1GBcORcEdOVGKPbJG75dLZX8fYzaXKYUbS9pCtAzU3dYRMeOIKPqo8NMFv3RU0/kGQpSawLy
qPf0jyu/W5AFfxNKNHhc8/Rt3pwF7bNTR6CtkiWsjszPfEGI52K+DVbqHnUfFwikY5ce5aCrW7jo
ujLVDXY2SdPBE5J/xHz3jzMJCpz4prwY3iU+AeZfiulADDA5uiezmWATR+D4so7GjLVWPg4XRFs8
HpPvJaxfupoHR74bVbNeN1qfiYAHYpl5GCfw/YwgG8i07HaRA01hmHeQ85C/QN0gU/xjHGLJXOv9
4g8qaOEHxXsX3iTzckNSafMbVK/wi/6l/6ELTlHaBYLmyUV+CkgxuJjfSAwV8eeQJ7qVPK1QjzEx
nOR3ia/FwsM+WJaO47BNnj94xRNZgqcQ3weom2AO/ulSIaRlXDLOJ7ddq76EQBa2zFW51lJrdTbQ
XqGYWCjowgVp5+BtLwKpYmeqGurBADCtzDGoOiIVtjMrzkVvY5AJQgeXfeiB3iUws012Nih6PNu6
TNpfXFAP8dwBZPgjG/xKah163cxt5YVTpv3Z2xLJrLGS4ZnT9ME2pKKFupbJMxgwOI69LBWFhxe0
c8S8Je2Gido/DKrU1sKpVbpYBq1rily4ePKFZqJ7TdJ6MMw+PW+jhxDTaLV+mvt8q5I4cq6hRVFL
QCBO8Ar7JsKXV6TcOn4HM2/ogKt0tZFzTrd3nX10sG3LUBToT/7M/I130UCxpnZgi3o/C55c3WcV
qETC4CMXekRqPj81FyMPVtf4I1Vk+Qn2mZb9I5TAPaW7DF5d+FPSFxHepPmIKi8+OYZfQEj7+191
NQs1DH5fNk/vjQ+4tXf+Z+apTlpwxWZftuBV479I73e3hmnM6aRjmJgPvXQzaCv3IrGLPnZ4tZa3
VYJONcT9CvMNHraw3R4J6M+sbbOFIdCxi2Rn+f8+ExFPdeTuU2xCC9zwFwaYdvFbwouxHtIP/fqd
0sLPaCsvFdCcRSPeOg0HZGOXg8wAI602XYtyl3nPDHPV8ioF/f+HVHWDIQxFgYNq0+2ZTLBwQIxr
N6GPllc/L4ARrKCiNBAVkp0caYjfWojhsIsC5yaV18rqGovZwRWxZJ5s0HZN6y8pSXqBcCXZlAYS
GpROwYWGBBuyN0Tg7EgQU0vxiap1FZGS6qH+oy80o2ypmhcCm6r4YfD2Yr7np/ia2Bj25VoVknoG
p/wXf+lnJ8LwYVfGjZJQB5PDj+mm+29WmqpvQ1QmaN8z2XZDGbfCU2Gfu6JXWztU3L8Ah/CtuCui
oESzJu2ivgEwz616ABt2eVH1wdbGA7jlx2m+RUq+REWEyUnmntD3vfecs0bzgXYX7TZKiZorHsTF
k6foGUllLJY8GB0MQNCYaGbddbdaTj5MLWrifwpfNmqXJAgoqwRUNcnznGOp6tO7yMvmm3w1Db84
dXGnbSDlCcQ7dxi4GBgBn258VtOcrQPzhFWwUTQ/bmd91cY7WrljYd3ETRa/tY6pmXgLu6utW6pe
Y48Og1dVTvPh5xWAzSAtVsksCrhL1vZHO6HV/IiF7FTvMLX1quiKepGKDIDnEN8OV1O7lKqea2Q5
CnmLl87HeGDcPuK6xrtWNW8qcb9HQEjHi/7yFMMWAVk/6SvClKaTFa97jVeVJjCe6/HfmLtcLAau
YO2lnfWURYlWtmOCq05xwXawnFGzUdIUL/1PElXMdfO4OgIHfeqNo/lwO35QAA+zu9bBrJ3jz42U
m+iORAIrivh5QauRJQ8AnXSmTi7i2bU0YWtsEVTgIHUQRFO5hW5fp0KM1A9RDalzW7qHK8kvBwEP
kVeV80FMyHsF9z0k5tJ/5IwXZp0jtJnjMRhYUUT/w4ReSHmS6eujwq+dFRiHC3Ncv6zqBzkgRw5h
MAE378KLJYcbHyZtRe6uHrkAK2KJ4uZvZvArcDKWNU9egzPWwaf3EzZy1vRYFtigpMdro5LJSgpE
u6RmNZSv/q40JDo0GMeU13mu2OE0PhUqPIuVd+kt5vvdIzza5i1wGLybPDTXYDh4QByAl/ycpe9O
jMjvjD4baFXbwCO++xhKbaXev9qfQKLoV6uZ1/BOsACdAyq6jQVRfxP+fbicS6QaF7oJt27wXT9v
6tgRJwTZaM6aWwjmlK1IgfXvcgTBrrq5to98MHHNAvpf+Jer0JU3VkeIPFWI/CuX9DdtsRwrU+AI
VLM+xcngbmw5i8WSUpwKsc9v3SNAC5Dw+44kA90Kx7zZEPHTPpatl3y4AzVQQUt+vO88QO+DXRKX
KDjiKhKEEEGJWcWWzX2f9w1RlXvV95SFSu5lrRUcwK5ueTyv242fAuC9T0bhzm7Y3SngWDxLX3Pv
95NwIV73Ao41CCFA0So7mC+aDaUg7tGGSi5VxHeVJgiU0ubWKdq63bLx/Mixr1QOcVjvIec9G7ia
lG+SU2YqqkDJ7p6NjMaP5LT07Pfr3JlNL0QtbLnkUK/YfpuNZHCyJf4Q4c2qt+qKxVEaQ7wTu8fC
+KWI5ggO8/8l3Skkw2NLHuWuEh5cYl/DqIshLA+HmIEG87cUEvoAxNaWAO79/F4uTUaoWxH7/dix
dcNqBBAE9sY3ht959bSkTqmMKOA34ZRZMhCevculU3zk4N4jtQsHacZh+CYBt/4ta1r3lxSPmQcU
uft1pDnP3wsI2TH92D9OVF6ALTW+FfyNUIUJ3Kq3oZ40zqulTNiivcvfaRtGGVSTFGqhxXZsK9tp
YPZEfmwWRu57tHWISQL2CCMk5gsA0LASk6IcKOMcLK196NgRDcSXB11qcTF6rXvAXIqGv1Kr3AjM
KB4HMilN1crocKQ0/ad7ZDb/2APq8Dwlv21kRQ/mRtLPMk58oY8NxKg0E0L585+WNZxn8hPLThBy
b97lhVz0Qoy497qNygenHqxx4XwtiOAwcWmJ+NBwZzWU78Smawq/3Z7V9xZ4whRMpiTCfu+AKRfK
EUyLA0SnvHtzmOPRp2p6FadFPtK2Jtf/B0TfK7ITKKmDIxEF0yRjduJpbPcdlB9l2/M4YYb9NRYY
s+ekazYeOu92aLfiaEBCymqmMQO+sgZElrbOE8pgWYRgpn7sEFdL4pmxn79C6xvP3cUQsH6Okw52
UfGpx0FTjDddagixOZDHS3yI7Q1L7X3VcaSdQRkl+gNAf5wBSW33UfkCuJkDTC0BcpyJdjV/GB3U
2WxKOB1aFCB7kM3ffEvalcVgAloPdq3CjxEXQQxID25KEvnspjRo8ZNCdedT0Ux8ciNFMqEMDItz
oDVixIfm1fkyBmBhydHxzZQw5gfNJQSCfcnnjZxTWYHX3d9CVLUJREaEM7AP9Fx/8PP3QKj6gR93
bvyH413R96Ry9d80G2ove4Bu00J7vbG36mzdpUkpMOpf3a7CmicAhdc2q+P/hWe++255/ZXxKcE9
7Lp8lOnmUhwmsm86b8VBIDsLolyl4pDtK3ZC+RWCXPXC3tezwBDF9s9t2Ku41JmRzD8Ph7vTnKC/
EsLkKZpBWh/80ezFFd18AQXurgaW/ytggX6rXPZzDFQqagpujWX2YGiFkw4sztDotCcX6Kd4n4jO
l6olse4s2j2eB6+OHEAvGAkLHQaHB9kbxpGQPXdpfYGJpix1VMHYHxaRzbh95lJdo/PID/n+WMPy
+5GZwuVsMR/0p/3zH42d8ba+ouBQAFffyYKilRtzHxTkQeH8bsA1PyLKXaT23Y45nFxPh2dkUaWa
fmWFJbJsgMeqeTIrblrPkcZRqU0u2H9z+P/O81J7EHRFIqZFE+9mRNUd1mkNgXWII8x5r23NFnjo
6urWCTIxzL0/8xiHdWQtyGZlo0NLHtd4d2YMBmjpwgRTEZ7m7e1WfN0HTT3q8xNEk1vOiqjzeAsq
3xxxdjwXxjJUWIO4tZyo5If4vq88cpDI1+7pMs9XYbwP1T/1iEDZS8d48/barYvOyxCPyP4Sf0vJ
YslZSM/sFRHjU72npJ8zm4rVNXlID+B5yUXFy2gaxUnlc82r5s/Gw5BZJeAsxK08UvP968mlfv9F
KVSAokI0ik/6J6DHfMwev46pWzSpOI5DJ2TylkHAgAB7m/uEUt1ihFlNodfb4onDrjLmVNT2Ag7I
V7t1TeK8wL+GxlmDWuDVA3uWTqarFZksmqd7liofgUFApEzrIyP5NhaksPaXp09qXCGth9yVP0rq
vUpUTyAM2BUUNVgCjBtJrGawBTQOFdaeXFaGDmIAnNomU41jj5n/PX5HdjN/I8vgHVDu4vaC2tcd
NiItteLPFMeXBKxj+TDi3ufq6VwHxxnqv1S0EiWbXuoNxkwNAEEZxtnfeXTw1MtfEiiT6xQYnKhQ
HmcF4+0bJ6WL1RWi8MVXfT0z+pzytVm8sQ5+OeisDqAGhKpuJudMNDOpeY/STSs0RCaxDe8eYZAb
UAfgBCFiWZsQGwhFBNMMinjI9T7OKMqa+TWl52ugwHQ9eXSIS67VdkU8NOqCkMdc/SgqMiDtWXuI
I/niP4KOIhRH0v0BAGGJJ6DY1xXWddjdPpMn5gtk5DMgT45ILZJ3dZsierFrJiucjiQna854qKbz
8tzWIt3s4vk3aYGKHTgea5d54bXBls7IzVVxuZ2/ldWfKYXTG8JEsEkxgCu9RNiqQ21ed+wQk0fU
40sp5MQ5drJm4A3j13f1MET2HuzMy+KSJw00u2W9w+9z8a+GfSFeLLgW6sbyxQ7dWa8FbnpjbFcf
/sAV7Ga8coI0TiH8VKyzjMjoAqkeR5LKBnlijq5RekrR7ZpLUclCrQVGtAzO+smIRLuYVXowBjwq
HohO5jpSrBwZYP8Xn6fN8/bpjANS6tqTTtB1bP3Qpfvaxt9ThvBDRBFkwi4OIFoHs16Z8Y6oLIkr
q3obNwHou2qWXrOFJcgC/ppeJkZTjRa6BsIa0+7jAYaGYGYZivd50hANPkfENSK2tD+B0t1ZH0k8
a3Und3F1fpNgwdZ3xs9lM2lpceDYW3bgdluQ+bwvjYQ+XJXcR18oZjSETgRxMq/fjJHh8vHw2g+d
ozwyW67DcXKCiTOIiUqVkK+hW/JyN9RDakfMHRXllQQDlpVd2xNkPx/eomZXWkTrMKPucHB34N34
Bvm4mVEfGvB9eiKFF2fSZi4WSzzbSNoMn1VBhRzmI2fXH9/ZOQQiBjVJrJ//p7IS4iRqGfXbO1oI
uZzEe0PPpM6yz3atNcFj7Ce4/qH8iFDqyQltCjSRfQEEkMMr4Fo0nNNHbwLJpKBLE/IrJ2j94kLB
c8Hnm86mPeh/G1wEXJuC5Z7ru6RD9O6Danl2pQHQQhibgXJRIkDTjwRSK+vY8+VeBPFPBLO3hiHe
tqCbqDstNuIpMdxSmE13zFWR/TNpgyrADL0MW6/VXFEy9R4FZ9GaEMB+UnCsT6s80IIVCClo8KZu
ILn92Vjlryk5JJ76TuZP43NR4YXfrTYV7M9LejuV4JbZZqE4sxAWYD4F4s9R8zxFNkXoS1rApEMl
UW/y6b0Se+I+D+J7CSAjZqDsJqYWMb5BCRaT9ClP+zM183SLhQ+a48bttx8ypgOz3dOZGL8Rx78e
aUgw6AwROE6U/i0IL+G3vqHhQ8qxz7GoeYy5qUzDg0bin2ZvBv8BwgJIdCxziIwRTsVb5nrZTmjQ
RCB0WKUV0NRBthLuwEhBjxPPW45KlR82atrXi2ujlkMbSt9Z0jByHVVlJegH+5PmKLe3VLDQEqjc
0Dnj1hgzwlNpmBMkEflDlOZ1f6u5CS4jgboHrm7fypoM3Gzy+noxbYnk14DQUJyRQENETHl33wjP
b2QBjsYY7OpOg8AH9qWCR09CoQPMZkGzJNF8jyVCf9UK91409TP9eKxMig4ktdxa2T5Rn5mkWbYw
wsIuDnt6k/cDrGeD1dGyboovWuYjKppLPC5moaFt2+xfYDsgMXhyQYxETBE7DTbbnsibihLji3yU
PelO4mVVp6akkz8+Ejt28SqBLf3bFuIz1GexCZJo1pOYO9kiiDmFfN3QIUM0BDVXL8dm8MRfk4Lg
62p8MGbCV8+Q/czbca7VAxwLUmIjQeDHS4emhuHZB4GL49LoNuCSqTRc0ia/aGQQ/EXLDPihMknQ
0D9U9xHan+f3Inwot+npze7gTN+nPA7wTr/ofhsmgci36IAbQc8zqyl6mIuK4cEYDH5QLTwPEtH8
gUUpYDv00HSCWIgM2pKoHiuj2CUgFi16EDI5BEIwFzM2vHOQhoJoFyA5QTZtAclgJV3mqQmSJ+Al
FqVJXmFw0bcR/rxkF/0ioV8MYIDZ2Vbh3+SpkV0a8xbnUpHeJDb81FdubJA3W2d1K0ZrM7Ql4gWw
EC5zHOsdrqaCnIu/dQ/TJsEM0EnYp9eh++q+kGY8f82dtQNvrEM9fgbJFJbUN87xhykF4MGdnr9D
PvgYZVFQLbSyZ7z2gutNpEsv3NsuSQtL1ZRdDWTzdVxysOveMwTF+C+tLgCU9YlZkj5092Nq54E4
jtHmEj4bQQAlaBTyhTl3G0oJEJutK222s9E5W9z7RyUgTPmu0nxUvT+MswMLbBVajywWGWzWXnkV
ccZ113tp2vNv5OAD7ln3uWOU4USpTT+pk5jlOblpIAfeWVjAa5ZEsz4DE91OdQeqXF4YXc5BnPUe
cLiQHVHTlW4KnWlMiJRuNWrzlYQLBgbFTTT8OwBEiMGIVDE59+Nf7Cflg8ZnWG/p7GPAUP0YmSPV
UOnKeEJhF9W2m+eEHeH80BLYL+dFjr8N46X4JNkU6JjCfAc6Q7X/O2sk8Y0zBC1lFvxxPRLgCG5B
p652vQPv3lCMje9E4sSjfmXLTMO2eWK+kbhY0JT96DB87wyoipf9UOxn7DZ/ueDkBc3nqkOIQ8Pf
bCMkx4GH1du3n+E57kEtoh/DaxuypuzDu4LLStk2faBuYwmwktg60HVErwD4DABl265uoc9dJht+
nQ8fS6L0quFezz1fZYIUG/V+/GMCGZnyBFPVqI4sApdLxdusPuS4r4qKlQqu6yXBHBIuulBr5pzx
ISWhbhSo0sDFv6BKMaLcc34HAxGP9fV7m3zGc/UPvNpTAaeZyLUd84chPh2KUHpWcJebnQwi/6iu
W1OrOwjwO3H/hGsFcTAecZ4+kskTfLAA64hfLMVkykokrGgO9+AzvfJffOqRbTArF4IN7/u2hFUV
2/FlH71U79+9vvezOnWR+eQYK9vJy7XKRQVKpWsE+q2HlZ+CCX//S7J4mpogyqxwj1dopBPPjxfq
R8RASHpTEn/P55TXj/RittfzPn4P+tKm8wlHKDviTiCpR2eFUxl5AqLr7/M3R0ajnYy9q4Wz9yMR
nXfPBMV+OflUw0EudtjWOumvbxwYfrcCbrkcdSrTCSjmOV1M6RNZl7gAaWr9PtXk1rHRRBrdO2uD
AMk4tciIRsr7bCUc3DXLzpSNpe9wikC1OTb4Bqqla67qbP+1P3zBxjBhxncNqo5/BeeUf6p4F/BV
fD3ZQ3ssLjJ9IQ5q+lY7LWvRXUS5c/xOVVVuXc2xTKpGPo+9Hn15OOf9uAkEqMCsd+QpcOOEfs6X
Ed2JW8x8qdApd06PmH0CoKG1TpsZyyY9hme3GrbfeKl6WuJJqUDQJ7Hx0xA5P15cyR9LMFeC2qM6
xRaV5x3h5F+1W0Ptv7Wvyf3v+OYvCoBRx43l16SZ+xeEggUaBBXc3tybTiNSChaIiZuUd37OI98T
aMjSMzxNTNzmGaTCoW0SzLmx7P/fZhOVfS7X8rh18go/aozbYRTLTqk7uyjdA7C58QeVpvZpAjsV
DZXcOEYX9K5uhcTha4usUvvRUI7z69SFDbwGeR2wQCkA2hsQ64onRSxzRGjuJsfezyPXvHGrnYhz
WujSNMMzxAI9dh++E0997S31h94H8YPbJREpMyjScIApCbqyejjiVvjcjpNR4wJjDvE8HQ8W4HGI
HpvrrZradxqXqF5M9hmSICSejdv4VmRHAj/6POIZW/vHMUmM2B0uXITCvIzUXCMzufe5WBQ4hERH
kzJikipYBswlWj/F7xwGAv5QGl/j8OPV5XUtri+hRA6n+ZvQZOW81Dy7MX/fZe20I8nEXUpWo3Nn
FjWOYKZaLTec8ToCV3B3hATeJQPY9mKuC1DWWveoDrWUO+xFyTbI8Nb+e7/05uT/mXJAMxYxJ4to
HRwjeOl7m3WmOYYMYN5/v0ZQ8IiTtfSvSTmaZtQATHeblezslyRMkYx9hRwPuSI/MveoTGACxy3g
QwpieIpDgzUZnqeA/2PSvBB90cYWpEo8a19MT27xT/xHPNS2dOKQ8DChzpAWo7Qj+PUU8Bk7UanP
Xu4pLhaNnGxE34GEPvNXkV+kJ7+sJaQ3OEvL7OFmgnkDb7vspNtRy2wtZbrG8c1ybqXzw0Xvj9tr
Gp29b42mdUQ+04VJA7c5BPMVpf7XmWZht/0NGu/wfrWPHZaNWy9DFetYzVoFVxzF0EUdJsOn8AWv
/LFzDqPg2AU7QwEVUd2pe0xBBZKOslcljSCL1+RhmRDzW5y/izn5F09cRFusiztdlx341hB6SJ3H
2P5XYBoe4JbByeLhE90uWpyuM/Y30QG6IZWEuR6cEXCskrvfjjsD/7+Be6Q8ngJP8qwhvZVRoKV/
sbHBYMb4f7vdoHsxg32K8aR12Qe/VAwM+8QViS/wEOXGHOFAh4cfUEJia4GN+UCkINifKaXDXCaK
AO4EUr+Ex3q3f+DPPf/LVDXnBqYX3LPX4t1wWpK1oVW+3X3Ax0OvhM3W/ZJ2JUTTrCehib1Kmpq0
tBUX+xQjJzjBZRRj76PIPYlhZ1g/8NSiL6iMRkekeCMY8hJv/0clEOGg8k7sxhq3GpGQ23GGAc3A
cOpnmtmPFOQvAmWD0RAVsNmddUISEIAwrEOjMzOB22vjMXgXDK4G44O2uwUzTp0OAN8VNSWGD54d
o9vJ9QOSNG7Lc5hEUG3x3nCGg2aFSCSO20vEI//y4KFyQUC6/ek8rCMySEgewGQmLP6YVBhCXNXM
QVPEphphJt13WqSjfvR2tnIBM8otMBvztGH1kvl1kJeaPiWYYnop83fsBIYkrVhj/rYiXZgdhQLI
FWC2ppiPhquAn5t5PYPmzljKGwDsDryDl1JSU2JxTcMfnmzyy5YOWa1OELxBT9bpV2it2O7nAXtw
WOTmDQRJvSGxboPPGl3t7Qz52QVUmRU6s5p5hNmb5js2NDT8R+EMpmPJdcYVK8VIbf3MpRjGe+oK
IhZRvXMQ4Fs3S+uxQC2XAIedYDRAZ67IflYjAUpEhyoroC7COMtwya0jOr8vlnMwKl2zI2rZWUyM
geTryPWb5dpcKZHPZTDFEs9734BmrqGhMB7i99DVQZKM6unXvH/wIaVTHkcc4mkuomLlJFvREwBA
2FIHwxDSUx+tQTg+Dhv1xLls9yUg7BeFKH7/4UbEAH9IgD+iS65ybvh6kvB0DAqUaF8ymr2ItxVK
vncgOksC2KkpbNEu/IwGtMK5exge5CH9TPtpVC+U/ERNSWthIu7/v8z3bHAxP5jT/5bKUlajpSsn
rbfkhXh5mcDX/is+OamGtgXaXztFJhKqOo8cZMKpWHODIToSRvjW3E1iYadYwaFrP/ULTh4IorAr
Z7u2a53DtSMcMFjcqm0cDxT9AP9bjYz/nTmFdFMDxQOfdxMKRfZZ19zDewucFnttA0JcYsig0ere
eBm+F+7u2gMdAB5ezOeC1jUKC/GpipWMRKUVmKIoyEvNLRJGW17ZdE7iJQERsRb2653qbBs4O/Iu
aptvoxabJzD2851oFiMDnDDuoNYxPAHvKY3j1hGYoR4IISPU6iqNlbj6XLpu0+3XkJdkzM40Pfh5
M0aPjChWK1m5lzVz3kq2GapklNBNkSU1lhbYCCrS8ysRsVfQysYivAqbuy4JNHb4w8vXFNhtvW+J
NMK43pahX/+3fkczGBRwKiUMNWsj5HlQ+1ao7CUi/wyK8UZkrIAVvWmlau20brTODYpeDQQIfxZY
o5JfiH/jwJSab54vTdH0yWSYbwpV6ORWk1gSHIXyh39qW9+88I9oSVU7zMTop0o8SGYwA4YHaxdm
W4XMtl2NaVW87ODfsrIed8UcwlxVlndxy2a3uYdyZ2ow9H1t1HFaUDsNhO0VAyUa3S3l9KvERjeI
Kw/MEEcNihya+AeXRPf5/m+RBgmFUdcJfFAQxEYUHxQOPnb+dhvHQLSaVrXC91ORlNYxAg4BBNDe
ZUqR1bjAXffiZZjZtx3VFH3xHNi4N4NrP7N1oZwMh6+L+TWu9w0ArVKTk27wG9eIh+7DdQs8DXD5
MQaP09+VpxPKTU4BjEvxNHC+1AYu8Rog1ZxTwUVWiPQN1q2J+3Ns3c6UJbaHxtWLZKh1e91jNaVg
/Gy+xOnli4qzMfejfiby9zQdTxsdC3qejkCIGVxRRWAmoj8zPLbwe9aVXwgv0wHzYVngNlqs9xxp
YkSXDoHyG5E8YlaycsYGcfKkWfebFiafN0mSqAwEm9f6mo9/XlVtB2qYXxn+/uQER0slNiZGnoaD
u42VA3V7sttuqo2ZQrlErCLMHLBPIcDO6/Ot02YyqpMy55ZH58I8aDXjxFgj4pEqD2XhHq5oF9pf
5GihcE6QWxgG75o7Q/LWT0UhbQMN7Yzttt0yW6SPa8GkXwrN6xKYX4vR3WB50h17NOZxUz8VUKjg
f9C+7wtPq9bc6YnNf9PF/qVGP73rCAvAVxaICwyVy+AQ+PKklQTihHIxCsZKZvOgbmXiz+TtMM4q
vSU5qkaWxkFFGtCRseHqCkpxUsZmBLkW1pLeFlDlck8sB8Js8MSlhex5E+/gnQKDccsipiltbdAh
cHX9Eh1xSF9d+whWhjRlTJwSYb3JQGgm/KvkeX7oHHaNjst/iuXtHSlEoF+CgPQF/9nXeWRAGoCv
fJ7MzVkT0B7q4z93behXTVFNZPPBMBocPwykdgNWn9/Nxeb1Gtm6b9CwvYxWXUYD8pW/xflf8ihY
apq7Z1Ia1EaY1v5t+hXmdk8sKWQgYLIrZhxjzIELzpJAa/Qc8J7PmMvjYOdVIsexPEdpnII2kSRZ
3dFebfDuq6u1JqKXNWTwWifVeTs2aU/J3g0yqtQ8WhqfTfM/zOzYjOYdNmZzqb7lSU17iH/3l6oc
+bfD8XLmiAElLKy7BM6kqSLo96Sc/xu/TDHcliCFMATXv4zFArRKkf6vCy9lG7ByZAoU+5BjjKX6
CrchuH7iVmk8u5Fr4Eprc/TK2VfxoUORRvcnKcd99yHerN82m1qLFtMnDP9J1xxsXVjC3Uo67O5B
CHProvHsCBcCvLVtxW6tnlKDbzvVm07YFvhT/L8DwtSexdqtvB4S5jXXtPZcNH2QcKE977fw9w4y
8G2E2QtnpPsnJliisQr5EGgfqoiXMJDQxoMfijNM1QQ2ied7yVeCoj8of6K1Eb+gst4FAVHCYgXH
fMfqDX1KLsx9yWHtR491BHhjxVEcVNBHke1xKeBHSsM/XKmEnCtQWapWBzxLo0UQMI+sLGocrfvB
9zMloNh84GWFmSj/2dCZjLu5RswsTf6Mrfi4+FVGGE2s/H6tbujStBaOXJrgnuuSGeF6SBCGbDPt
QNdrNuiFOPEFOptG5cylx+iRhxJN9ZKHoDLQTZZQ4rokeW/tBM8n+OD6bnsfS3o3dfvaTQfEg9qz
yyxrBe7wJWBrJpK6xD/+oJ3LWFafVqy0idz1V1KfPfW8ESjbj8Lh/z0SFMEBWHZOxZh4BVc1tvgs
QA5h4EgPqAhvJo7qscitFjA5qWkjwZ1SfHNrojbllTBb1/hihlNDqTTNIdoeCKr9ZB6jkSqmYe2D
jUSVFf/WBwX1iJF10CQrUZKNCLv3wbmZ8e0/cWPNeaTRu22UJf1Gxu4jgtRjz1OuPN6A3zDNlVV6
M6TtFURbYs23afRvwswmpRs17Wfxw5QWpr5DE5oi4bhk4mZPhPqt3qcTbxQ2HF2+3V/cXcx9WrPj
H7JAT2ccgAftyI2GxFNzIE8u/uBkNULtQErrLcHX1NbtFMwEVbVyx+EvoUYox/KGPSbPfjGVLCs/
8ThZY2BpBnR38m9rgtB8R7nvw70BiB12mbpG5zt0525awfNoi0YC5V0FpKY10W9nVK/v8Tgz8qof
KZG8uL2FEk/XgJeTdwfl+R79ZBQnsI5rdNaol0KCuLcX20qtbUALxQ50LXRgi82anlP1B8kTST9e
aab5cEE+A1Weaherdv7DcnxzgpflnlUZuzWTEzpGGjevYUbT5THbZ8MYlgFm5LF7uRCxACO0Wb4+
OfERafiu3ZPDDkd/ccb4RpjfJsfHY94dWb88KVFOMdgSsNjd2LopkFGLodzjPr4ass89cpz6XX6H
Oa08O4tlEF0lFQ6dZ90t/FK7SifYKoueVY0cEFmOY4C7UQ+eaPLOpPYeh+WG/SydOpQhU1OFmX7S
BPDGJKI6xA3A+n3ucTLmMFUzrSkoKZ19DUbOM1igWJGjulOZnXtK3SiKzZfTkEWQTB/lO4/bLW9c
MwqwxreugITGcM+U9D+0sx6kj5S9Or3ruZl9ZMDPMJ0UG9f0FjQWLu02L6Mi3jf0G7v0fusItkkn
kXGh8T4vW9u7lbW5Ig3MSp1F3wluZL/6HUAwx1a8NE8iXLlhLEphA9WXyYq9TP2qOQC8yEzKoxjX
bzntpW3wmpcuEyd5txLO2YbD9JMPLjSJDD7EVxRF3yvf6uhW9byyDzGJW6mXif2RTieoIAVyIYhW
tBgLavySZgLNWmo1hBq6fJ5DX4pFj+UMIgxIGqky0NANu5VA+6rFYW6h1uY58B5LHaMJTMENHyGj
xso1iLcDstMseQ9UN6/AZJOEBpWitS7rcJUOKu2vBwvsPQLwhtMHFNAHezU6x4ENyvVG+MhTjgeR
obGUn54/o7a9kV3jclPCJL7ZibA+kMTw8bBf6QtFU/U1OpKAa2hkz4Ct5sK1s5jAXJhBBWfQcnWK
32Egmv/hfFjeSQTzrdFEx5SsTNxr2lXQTLz5UomcxhqjI8g9OzN0Heg4hfRN+WY5Y/4yP/IfCi/7
ZlTIr9yiL5INO9lVZZeSEyBf1gSCWLLX85C//pTrvQ02Rewxwe7sFDpC6G/TJ1DvQmzEdqSRF5lB
MXtPbS7e+JjC5PephS1HPYlhVEgj+ONbs3Pfad0lq6F5cOhDajjprvuRGxjYpAllcQQ0AvzFY9qN
mpnbFN0HfwcyQlr1eA1pS204u4mNxNYzXl9ZvOOwNCaSZM7+C6XisWwYQ/s5y+K5w+1hz8+TBpQ3
Aexelw3d5IDw2gUtIgw51I0/ghJHvDmLyS2nOJWXdhT9tqvrYjH3x/SH/aXkJO3sFG+H4FgiNluJ
sOWABhQdfSSyHE9Hlj4FGjbZ+yTOFEMCfBZzevqvbSpGeOyh86OyNLq06C6gYS7rSDMnimJ9qB2l
l8dCwGIBkoukcw4s/MW3h6/lGsdLB4gYhiWYYbOaYQ9DeI9Q2nXxWsQfx7Puk/YVHO6iNOi1n/iO
iP9R8oN2N5+3RHmgABeUxwEY0Ls0YzKhqxCiX+e8LQPx+XOaINUF+a7E4Bcfj8M2V3H0U8nrwo1Z
snChRteU+ZR6l23zHUq/WWQw/GJtWuD+vNYyyBCA71Acl59rX2UezFXt1U4k4QrhsD3dbOEw/4pO
wdf8cvAokIZoG5W7LYX48oEYY8QJZZrqxsHEroTiIWFmx7jFfr5BJumB/IXyc916Dwdb7qlOjwjr
1YYuloUV3FPCcm5UcQUdcmV5ORs9VEGC2WirPCHXQVBBLKDX2Yyb7PJdujxwxzYYN9kf8QNeWjvt
deqdl3jvOjDy0CIsrLpcqG7mU3v/3d+qhQODGTO4T88NzBiM1aJUYvV8QrtXBEn6PKQJ0oY0tmu5
kUc38cJIaRRmKm4MAzYSQ2fn3wvJzKss/iqvont/xaOkxlw84A3MQ3iRPrTsyCH2LncbNhYt9wzh
Nr+0UJN3Um/JfRkdysI+udiF1IQfuaIDyzeA9WfsvVcHUyA0RgG7xauaJtIjtzBdWOP4GysQp5mB
UEqKvn3AQCInO6zw4I1A5SLAGlZtd3oyyoSPFOCtOADi5fbdFD5AerM7Hm9cINSOZd65HTl9aD4v
zcZoFBKcZAijjzuvjjp/qaCe/2QAy5+/OtWlFXqilxIK8qD+/LBs2oxAp4Asj9ns2yFSIKfqDQCz
GdGcq2rHIbOW4NG/aRviT2S5fY12PpYwYdrNYsOQQ140xiGeSethZBNEeK+8O5DegIMJ/lS9GINn
FCoysmuq7uhamYRosINdeYX+bjCgIzN4YGf+9VlKOoyyB1NC2D58tk1814062cR4jU+uSO31wK6s
mHKUtl9GiGMNs0brCVQuYEHIT61ntRpbadLbZbizv5MutTU/UAdzRRdLuSckh3/bp8ylX/LpThnI
FAjX0oSOhmCsCdC31ZB5W5ZyWlHxgZidHzLcv3Eg2lu7RWGxU4FrDEFVx/bruD6p+LLNHr9KhvSp
sKPORSPsAYxoHwr0ZRmshyMs+3nmuOsvKhHliTgJqpKr1PXn+2ZMBaW2AzhcNWKxUo1noIGzJfzg
qJFI62wdex6SaqyUd2+N51P9XriWScOeznhnmEycE4r+KMVP08VxNimHhjJUftWET6fqfCxHCNZA
FtMX8tO/q71cz8VaSlp9AFZwxISMYfDUKaZI1UPZAackuqzNGNKeFLRaj72huAJSzHK8w5OT1Y01
1IBOvGuDYpYrBp6A/wQWynep+MHRuVEljAmh1WSL6zBT537WU0cd3amDJkYQ8y44KAadeILEn3v8
gehoiUTnSIMGiHq9zE6JJteoE7ZjhN9J4zPGHFjLXUHY/6xfvk5S/M4j4/nphJB2CFQxTcuUn/yo
M0hTc38UWGBWhJSx51rAEI7YKIcLWqcOBegYeakMDm4Vn1aYB7x3Baq2DcJnS2kPGoMsiZLkkIO8
i9Osgv5rUjGThaFCBHmwFMgVpUH3qjQws0ltlMB+RktISiza4NH05CAx535ZSUwvq2dwPQ+2EwR0
JbQmTZlulqoeCBAn0WE169RdMKv8Stfv7EOSKWoyzMfT6TCV+z7CjdmG6VRGGF8GnS0XcAMJ9Jyz
eAHwOpmoXmTmT1DZbD54lj7SQ1v+ZLWO3BdCcYjMKKNYY/DkjGtEfgBPjcecMPr5MxjUJgXnzAjk
3voVBOUlB7jroUdXuCdsJq9PFCcPqYQbfzkuT+a+ow9/xaIy5hg6qBzQw5JipSazJ9WigFbPPDg5
CnBSlIwlUhwW5cnW1v35SP3F032hsYZhr2yoIutJeJ9J8oKi0iAelxnRJ17iuldQVlABVQdVWJos
mwpcW7BH/dmJeoehndtfAA0CfRMWrCk2RpiRqfkNqN1ue51rkI1bi5ATUUeu5NythmyHGMmAC9K4
7xtC+Kae3s/r6DhBLQ8D/Zu8TWartBEg1srxQFUF708LhymVATU5gvysCzb403zE1KiAr4XFnDUE
ZhVQLlqe/w5A7F3hzrpMS4OQMP7d1+GOC3eDhYKHzGgk4in3ffO9363O2kukMxTKxYBvGY+H3WnM
5ZlHf4fTRRCRSs8XHHR9H0dDU0okdY8DCC2GcYuEV7yAWGVp/HOVjqWXGPxVakCN9revJHzxveBw
3ncNBgdkAxQDH0nPwonjYeKLrZn8PGv3Ulj8oJBjq6BK1evMG0ILwc/swF/dvlGP2lZtvPMG1n2p
RJSLLh3rW3NQwm/FacAEAAIKbOzDPxDKnTDlbMsi+Sftb1hvVM6ncoFEOJRwRkwe1KjftVN3WNzy
VT9nhXDVz5VKhRTYHEeDeqsRLfQil1Pj5O4aQFTEuWPzP2WmZeRSUCyir+KnuaLGrLGBXbTm9yNL
fmeXBAiKHBv44liTxqyVdvYabkyPdVNcVz5Z3cjeo4nfU4owMCC9MlkYD7lxNT2YpM+MjLmGu8yy
zDIX0+UeOrmVU/HewLOjBNp0+YiBbaFvg1FSQ1daa8Vo7DoFxGZtj+F//jU2/fAyxmu+/QJwKjrk
2EHhdVvI6qfM6wYaIoipzSeAh2F4Pr2+eUmW+pH4PMKxbLTm8Bps2e7kVnTjp1UxIyNkJBwLbh7G
ayQJWkyMGEBH9eWJ5tIdgcJis93fmxVeRZF8dJ30NpLY5rmZUQP6wgrFPidwsvVusWxTAbfyTHzE
8SPFhWuzcfsjCbAe4Vn19n/TcfF/nEsZFM9U/Ex3kU6YtpvNLzS9pBfEKjI/UkPSisdDC2XkH3f+
MEbQhIG+Ch8MZQqxTU1oeRQ0+rIIM7O55swzdB6kLuRzJWia1MDuUnIxuL9V2tVb/UI+ZZVnIGnl
6c0cEqWW8RSoNFhx3nCtCVcJnit29wSn/JnARpSaPnqrE9WYRBoDReEvZgqgmrocGOojUvYbFZXK
kQJ7xtdRtxlmZTnSttKg7LTY+0uV5biMtTzxGbc5+C7aOimRSRmCPzZWW2xv1BcoaYaEysjWluQt
eFgNWLaWpeOA1/mUHIkG2duhi0YIJ9FErwKinQKy+VXF8c0BQCuuFsSLcqTbupx+gpAceDbZ1sFZ
8E9r2w4Zn6NzM14ntVsYMNbNZ2vH47bjG2nIkh0heZbH6H6IQ329VgV+E6zilT1mG5TieRTMX+gw
/6FXSeEWvp6UCe2ffnU1v8zCk1y1rz2gKpUPuCg3ggwXO85Z2gKMiFv/YPD8rtxlcD1dl3ycXyHU
hWmpHsdMLLo93Cl8JwpuEeVtkM3TOl0BCwr068xm7vYBHZBEIkD1zRTUewolLGp99vpGaQjbmzl/
26EiKwxhLZVfogAmg9iIKfajWCJ3GHb+y1SzkXIadPddr2S71u7+0TyG+NFIdTrj0dDphraJKLU8
7/tiVFQKxx8e4DXrQT3emaHEgeXCdCOknr6pQnHZNpuJuXO3PHsiws0B1WFZEb9hqrexK0WVcJVS
BB7dBOa0UFiVjkpCtGgUedgVuGI2xUNpnoTsmQfwp7v2WiZxYZkWp0y1uLNHmcekBkt7wPY4j2Ah
WIR0KFzTi3RWggbdrZRjRi7KAnUOtGMT2gHnESsVvHzJ6RN3SSCQCVjDVENMIQmGBTYwpHcc6Ahl
3E1AQfEZlHfcKoOGApvWAE5nOagANMp+HU396pTxLL5AjdRYXm5kacCYsDnSgbtZ7NGcU2J4LXwz
da+JpriqCmOl36gNj6z2EbvSbKX6jVIJTDpFgawizBovAZcwmbD2TATIp4XZ5LazZcETAoK22Y/f
9Ude4U53eLUfeFdNwnvqVdD8Q2Rv4BuVc+LdbroeTHl+qQ/o1i5H73i6RBnZ0OfXN3kH5vK0h4uV
bM+N4nPawIayGjUVuAhAH11UYEI7M8/QUo/FB3D8g9ZGAR/Nz0+k6MNC606nDzKjRsOn4MhRoxM5
ljRswPXXn87RbD0gp8u2DFeDKBVXv3fEdaY5yMxy5vHV+pFbqZnVOJ68QHO8xGZuv7Jt86Pp8790
Gl5VDF/6ROU8/yFCSf3lZQt1YebGFmF75A398QqI0lfl4n+JwsLA95U88NUWfDrxHvJ6YBWdl8Qu
QI0DKfCnM4nHziaNCzrmoruxS/nobi8T3cgVacpbkkSHmYAYR7ygUytPDtIoQIODDBY0R1/mKI7t
XCC+N9mT4YxSrYh32AxttANrmH2DT7/MezSTz7DSqdKwBxKXgwm/PpZRmbYexrD1YBzBc45eOhlg
vDAz3PIw6NiYxoMiUKtyHTdrt8LtD47FnATBRCfxmR0ZlRNtXm1kwOOTlOHd9whyYps5TxQupndL
klbybwc2KsbxspQ3+fbE5YX7mFPZKzSuvFKww7nlE6VfgsNsU06TKTAXDXeJyYxCJnKqhNrCOZY7
BVEIjYWJLo+8LH+L2RMEMDQsguDDE/KrvlR+WPH/NFB59SRsqmxI6MHv70W5Hv9nxKq18PLBftP+
Z0THOaD5G7g//MU7xRfH9CWEIJMHe8a4j4ECRtuFf8j7pCdBwWvrEHA2XXQzpK9qNzygTbZWi9+i
xI8Ep4fF8MwdDX7u1Zzh+0sR3JALcpi+w5B/4cZ8NkITJHkQO7OpK4s9pNIsmrEZu3LByz6L3HAn
bMw6Nd4a1rJtGzdj3CsdPs97GSzplDeCBejidrKu8mg2wj9oGotH4GyMiwqOmPyLJfxrYD3pj7WP
EZJN8e90SPtqbe4catIi11TFk6v8HQAaiU+jkszQTl8wAYVdHovqVHsnvKefejKwBKpyn2ruJA9z
P7p08C1vbaXKoGPxozKoNMW7dt/uNYAQJjaqLr9StfKCZ9lQnMH+wakohHbCL857dCLJk1bEZ6OR
DDT0FkhPbxIi75+4Pyi2W8be7w9F1tVSlXHV9B0P1Y/UuMAaOueai7vd8Hsm4t/6+pTqu5vBVXmi
taHgOXmaFcF5YF0gzu4GrXchXOhn6KGEsEJcRhShuiXDCTeVXByXZ9Vw4G24u9zjayuOKi99hFSy
7lAlWvPxuy/hBZkV6YXxHfjUiPYnGVhEzKuqx1t3L0AfoWlkDv+N0gYppbw3228KFp0rh8zg65uk
coZj2WiSXhjq1uz69EpHWC5Q8AtaGgCrLI04DWglUNTP4GBFu/CmrnuZiRyoJ6r2l7emBwM2tnO9
oFSIfwNiHhwV+IGMro6DJs4sh50C1+5GOpwtNKvsTN/piDw3xSdG32l87pBp2E0ghZDIs1O1PUnD
6fA1bUuNfpL0R0XiuMxhbbIPZBxBTqwaONvXL3K2hmjIDjDEEHyjDhmJtcKyFFyduVbvK4n3fcJE
jch50ocBr1rdeHYNsO0nU+CSfEWWjA71M3F38/RXKqzzXMOn5Sm28zdNMdZGlW7hu02R4LYw9CMt
bnmVqWw5FYH3De0jzDBs+korHHzJKpMwPJAwLnguOxYAcULfjHNSFixpOkbpbMZNvn9dJ5Ul9GHI
+bjoLIYD0+1hrBKqNNqKBP5jVZmLM9miN3PXjNjcRYkh2Mc3AD1KPtRvtSYMEWEFY482/SffQ1Fj
NLg2vq/BH0+5QNddWiGkj0imgsPNgICZ3qGX7OUSyxDy0gkRML85twlc9VHeaIWdV3GQJX8IrEto
Z/63C4EdEpCZqzz2C/f8zeW+D38g+dP27ihr97G7T/EWaXLs/7itGSTxn1WGFEQmyuBOcG1S4All
h02NfGiyS9K8I4HkEVNoba3c17YaEikozEqRi5j5WVdlI1EbvHWk67NFN/nj84u53WlFiZm4audE
V3gv1+HOe2ZKYfhILBRgKWWtIA1bhHtx3cl4649UiyUf9DdUi+WYFCG7D0Cjy+1GyNWIuNuBZY3x
8Zh5JSCrn8JoYyJzjT6yDY01SoZpbPRIfZlhssdIURoof0z+XFs6uLc3kiH4CJ9uQ1gmN6R6dZrN
wVdFG0jUMuayfIvRf0ipzyT6J8S3rsfDx97/+D9FPQqGpNXRKsI++MZQ93oHFht5Iu0GaXsEEWJk
lrtX63lvfr2R1C6tkYMQ2nGCjQXe/se0FohUEZszfKXn+x+sowhDFVA9S2wKOHm0tgKXIaNFdFaQ
LmFYMhq82pBbBtu58jtRx89KGXOcKB74tA+SuA+2s7NkenXM/5NxgBh7h+vP37LpgP7aE3s7K2hw
7BAsXpYjJg2uXC2AYl54O+VZGMwjWNxVQd4ft8MFmqbx3ibCq89CqdM9lHxDs7yV4gFeohL75DQ/
VaZQ+TZtc9I5fpEeiwPh9KlYkpgMq/8xft1uCmZb4BSNnUwbt2M0VoByvgEeKjTUTYvdf+XQhNph
HFJoEdIiAcALTHKRT1FanlQNrepexC0403tj7XyRKVVWLjY4xOo1VipvysNsgwzXiAdd02HydJpB
v3d1Zw6rqlvpJsai1IsEABB+FIcOIgSIBwL4t6LvKNKdPLI6SmyswXbF9gLJIOozpWfLGbSaKZ13
qwJCH5U7kiv+cHOdD1a3Ncey2G8nnd78ZeRhulv/JPzHC0UTpK7jROXdJusVZ7dwEZd7Es1EPNKY
EcHLEst0CNAUXSieS+NuBTNZHE48o36IP+lb0rVduZILm9ngKT1qSorbLZlH4hhFfJdJGzEv2+OM
4cDhstJINrQhpAMZg74mp58K0NRO7migEjwaqP6+Ebh2NCs6TNT9FmhLdUCtxm5gTYEkLGxjfeQW
5zJVCmT5X13h6L9Fy4HL5/zWkUvXULXkhg7scSAK42ObaFlzrjY6aUZo61DGIZaiDjGnjfYFLPvh
kt5/coHwsGw2Sc5BRqEJaRux6x8RaJ1twZRbbNGNe4NWqMs21tf10ycSyfM6bJskQBjD81JLbc7R
0zYgW8QEjecwskuMQGTS0keUBslcODGZ0TvoSraZXToBWhBQwn+RpTyrwHvFD0yoZG7BpwYIzQ+H
Wth632f0AjzglftOb6TizPsU0GvIwglhizHAHMaCJ7LaV9eaD9/6VInE3Pfposn4ttiAQr1rdnXf
twrgaumsjFvtTCbNWh0MXVCODsHTx8MvU0Z2h4tTfPaOaXKA8LIkSgdi7nQJ30FOpES0ZyA4AvV1
xR5FyRcrX0ieqELrYbBE3lV6O9Q7jQWkS1fgcPXt5ykBJlYgt6S3vuF31fo/XhV4zYZ6jyHvh84E
5RdwWt1OjrSuupsjgbMuooomulJnuC0B58J3Kpu4BQIkLtlPlINqitqwTdPAmHOCYhZEApGgCaql
f8fjSAiVATyjjDO3NBv2eLNv5lUbPhF0vhJCBybPmwDTCVXm5tB5p+uodwVqYDsHaoqV4xddglU9
tfyl/hegEQZaIYH7Q8iVH5Kvqp/xyFuSkBO/BozPOESIDWucxFaIHmf9D6PO9xSZY0/717ePkET1
Pc1qpXfMHhIFIlKv02HZIdB8JwtMrth9zIsptus8hotWmtDUOOlNLeGevotfpwmEKO+E5xULtNfX
bPs7Ltb5JGTc4d9DNY2rnX+1RroYxi+fUUKYZDHDxhJwvYJLijqpqtsMyEAp3t6Bsd3sjbZjqWNn
VSaxj45rDUyH/7oBm8lE9Yex8jWOquZZ6AntP/lfnVE5B/vmTB8RAhuibCMosOx7b7QBX8dTpvFm
2sszQDlU/SYC7vaZq1CMeLAIJFHr5B7bROhWUwSPjYmL51xzApPNPoFQ3o8UXOwjILs8Q+xdTskk
GT4tAoHh+ReW+YrBu6U2VCanlbsdCInYj7zfdhSByYogehDTvXDi+TldEUlHPo51Qwhoxy0aeNoo
FhNA367VbNd5oU7qWpxrY7iOuhhlNSQzlgWIMESRFmlr2oAGu62MEHK3YzEnK4IGU4r8SiPmKr1E
weKBegcjgwIRIEBK6rxt68A68Wxzb9WXH8uKTQ112V3XCtYs5McZ82wQSMZPAM8SP1+IRJ8X8gqQ
drit4p+wAt1OwVe1NAeHpRd/PMA3a13aLa1E+ILFirpMqTqtgu/1Ihx7T/puFS23ZiVWYlh30VZs
CMapUKaLaS3vJWFtBbVSx36fK4EY7nsr+5HCf+9p8Gwp8xV8OgQg7CKj3eH93lHuNTd0g8Yt3jb1
sGFKg1bI8IRuofntUhHF7x68dsAh3E86rp8arURmmZnW2kwS1Gw6Cr/TldAxDqOLTAQaRMFU0tnR
flB/J4v40gRLcflxyNpwbI4QgkwBJ8l/PO4/eyRGSf41LniBrEGSLwO66TMoNWHPkVLTsJjajZgY
HSY/OIVl0vfb6j+mxpVBLZi9VmgcPLXP3pAXN4Q9LeFFTagTA0hHFjM3RK+wtxk7EAwaZPl17bWI
nYDTwREpSMfdSxfKrTh+IzUTded61jJUI9T4rxBsRIOL4Ssb+olbWEfLfjET2ddHRJCDU+pbkJaj
iDBdbBe5vLj8vWobboZobkgUTXnXlGCMrSE1q0priBqjCZLYauYseYcEqBEHdcZLXNDwGZOV43m3
kh74ijmdmCezibC2Qk5WJ0I9AAJmzxuKIgmwe4iHGNehu/9V3HKM0393vdboj/y6Icf1AX1GQFdJ
eSb/tzMtxSIylnjUIZGCj92HbO3/ulimi6uC5eLU/ROo0m8x/yL3La9pHNgkoIs0s3SDtUYDALnJ
a6Ild/11gfK8Io+FeNFcJYwekZ4D7YXGEcjWpty1OXGWumMZSJXQrbEjqquFYH5XjbMDzSPDV8sp
9scPLvKpV5efUNbeXxcse2JY9fwWGCCnPPue4rxZbFvLMas4+toWhqS8GPAp3FnvaABnPcOajlFC
SX6rb5AUYN7ouyZvMsF239VwBxiBW3xk0adAgkPiCUvcQYjtCZBKZ5Wj0JCxveoPVAiAB4EyR6BV
tNBEONrnFHHDLdO+mfucbKugi8eGORJiNsOAiVmsIal4gbNu+gLnvqdpOrno5f5G52/bggLxeCsz
/TWZ+5s0YOLah3C6UGwITjhgISMGCk+BhI5kgNuE/prJUL3iQ+X0dqo2JRms0xqABvD3pNCEjsEV
q7dOxsNYFTgdp7zhOvy/mOBGjYFTJKwmCw6hQWWEAq1MOTU2XAcMP8cUcaRebEU2b2lIerGgG/O0
tQbsbiQOANkDyndSqJtgeMuhgQLtmVEBtNhWQwSYOVAul0nXv4YdGp/nueu17smJVhkv7MGcTBIU
tpb8bobWaNhU2FDuPid3ALOtxQG8D9A3N40KlyFJ5XiZuaehtKGMK/vJaBxrnd/ex2LrRpqsvr0e
6hqX13jdakppbK2eqOvIdv/6yhRFDFbIdMmfFXC78wGGqnPmiIF02QmEcRSkpKvhT3UCmCPETPtf
YsXAzcemotBC/7qbI2VOXD9ed8ALDrtqcMbJK7+AWsczY3RWWv/s5qbWBuNkrU7bNUBJMsYPRTwA
GJAd4xtkObO3O+P2BrqoBUGLE4p3dqibMHdsXF/QeLCw8g3BIZ27gcz5OAAHsHeZ+LIWufS19+3o
Ht1M1+7z0zHRYT63HMbsmTg2I8hz6W1RJChA0IhX/mtZoX5Yn1FivztK2eXAK/D+su+WAvqFSJn7
D4yv03u/jYDbI1hFcMOg7aTF9s9tknK/XvHmP+iMtEQjLn3+C0kogzVsGNZ8vGxwmxcIKRP3uiQo
JzfkYC8d3zgOVNw3E4hKYxEf3E2XBkBJsU7g/UzWzV0q99Rsb/OWhMzLZ5lwY10gXQbRoC9XNkTW
iRX27XLjFoyFJijglOfnAJhIJrf3b01VdsbpGCc0KeeZGBzxEXQJ4FnriD1SzEp6y4Ne2+Dz8DEC
+9GfOwqhTFaOYROOvv7F1txvLTQ3Ojvc82XcNjIYkyFpNdNenOBiu9CDKPXPRzOA74mEF4Ik0EjD
IaeUpXqi/jmzTbdoazbGojiD5QHdLaIF2fvzCdk4lOtqt93Dspnpdv8J3XAC5U6w1CyEdzgqxyh/
NuQqj+Qz3H/lkVf6ZMnghtr7wztT6APaCeYLz6pXQRwcOhVoSxTwjl9KrzkhCtNEKn8sNzgM6QYD
qFeankLK7tDzX8iAlTfYDyOtk3QwJ8ngk7Dok07IK9DAR/QSImdEXI4vOARtpsdYxdvZHdD46IYZ
vaO7SX/uht1rQk7uCoPMrafDsnZSFTnk6fC3jh53XdgD7MNvfStxexhZLkSrmHgzJlbYEbpHUxR3
UK+7HOnGEa+gBtKa/xop1Qa8y3Ib0bLDHqQzhM+AvwBgN6DNWWxael93XJfdg+rnnDWlUfiEsb/V
aYe+XwQhFNb2apgrBvRSw0i75itS3L60sL9ufmtiJUraOC+IkQXpqKurj5LFelzNcjbvKDyz/6aH
mmVn7VYGsAxHzs0PYfe7UfXg+uymHaRx1guHHT0+nT+5VJq7w2hks0Vy+WROPfUa00ayOd+Df/yS
k/sFoDEs4ajMeUxZGhYbimLFJv4qRhu7pO9O1L4oPOWLkNezKqRTDc/B9vnPUF4YEr5hvE5t4Vq7
YmcocV6gABrtIQkC1+zN+ffwSNafjHb0hMjZxWhYOtSrD0g0FAOxOakmmSVVto1HEHamTaHBHm3/
UoAlXlwQ0IgELH0yNklUER6igm4qNXhbTF5c5NmgGIJ/VIalScF3ulFbzvbQhk/XFTmgi6r5eN47
LOsnEnaPq3qf6oVEl6ZM0WvJjDdKS6lI9hZQyRgvmN0oB/OgVHk9P6BO4tl+KQEs0uIvCcRwiUND
7xF/1pYOFxU3nWN7UakoiLMG4KnViP4YmRe+A1JV+yyZCObZ+eMS9AfXNhJ6JQ/ZNtVsrBDA+cpR
QV9/3yCwc2PRfse6L2rOzOYVrLDd9z9pJOXPqSmYFzQzr3DiZ2Twx6sr/4GW6yoLpRyp55q0SRmW
5w8wrPyYuMMOi5gS+2iIXl8hfvn381PlcmG6CFkZsSkmXp41R4UUCke5GOjdPanqwhGWDKGca3Mo
FSnTpBgCR63ay66+/gRDbxNfavM1rfaSf8K09bQIIw0p0qlvSwU2N54wSdLiGLcvbYxSI+FaU0GU
sdYV9qk52L1ZQZV9XrLnGWp+YaHHCVmTGO935UhgDcj6OySJ/5oJ9saVrYbGZY1tiKxdgIgGB+ue
F+kEGqPAM2rNW09m6arrUyVyTjUdAc9eGqe+ldKyh1MoTvO1xwpmTwINyid7AYf/sUgRXlBVSBxK
gcXHDLRzQV+YJ/xnUmRMMEXgHOzPEeF/Sk8GRfR8J3YuSp3oWbfLRsSCTs2981UpOzBqQZGVpIWk
g4EDPYn7+JQJvuFuT2E9g7fMYD7qwCpFARMlpxkNf101CES4pt/hdbP9pI2f7Xn17bM9XnvAVn4Q
B7SqH/CdtlLXBgkHAwEKZOdw2GofnZpP4V/FZ0DrCrft3xuC3YUgoITWJx4p+nse2cqw8svvrAOS
KWLDHgII6tAGrEwyvI6EMZhGx61kPhM2V1OZ1K9BrgFFVz64Ip8rbplryJWTlgNwH0sQLcZzJuje
ITMAjg/UUXligWAeOsOSoqUcHCJgTU48za70JIxko+ETUQAidPmteLR2zFs0M/Sxj1gDEJu3YKAt
3Am4xcfM+luYvW2nTltsnzVOUN2x7/iRmJo9HFYm30bpz8tLBYNBhV+aD9T7S40LcZF55d1itKiR
YUGT/A4nlgeJdfw/DAskzH/mbp52gkQ5nFPfvBrzMQIS78xsRQG08kJgmyj3R6kIVINe5MZMvoXW
glHB6IEInB3/OKfstWrIF7sxFOf9ZpCrLNGR9PZTxwIZHtsuN7GY9Tp9nnEY8ywxW1lQHTkwtg83
MZcV7c4VoQ9OX+O0hxxBUe6/PpliLUB7ogEzsHELV+K0VvxHPXHHY2h7UsA3BrTnyKQN7QWSVAd5
ODzdiDPEaa1J1F60GdvAqR9qDAj58T+J1XAI0foVStU8nxt3TinaA2WRpRYdlydwn4il0a7idd0e
kNUEdn07uDaXxjrzoU7QXLxkEN7YHV7EZcusmhUyP5elYGobtitYTuVfxRdvZ3zgpaLZBpWALoGp
pMHZle1FxrUhQ4e8m6KNFfwD7CSV0z0D08bnxp58aO/QbFPpaUC+BwFbjbcvJ1hQ5li5tAb+JFBx
cBAHOz/Y6doZXoGUt/fI5slwXRuoWOEN5bX4x8PW2qnlRKXJtiHkPQOgd5boOvfBXyRD1TAXYzSD
nv2J2pyUmw/9lM62KIDo2xA6W8jIcx4aHObKiwc5vMzpPDsu3fBT4vmdY+tndBkDJM4YrNPtqC2y
ofb662gPUOqyMGq6SNaq1WR4Wob+UvWL+98/wvhoiYS4goLok1H+QGCNVxSXEM83a/JlWf+jic5k
/vJoF1fAbquDQPSVoc3lDmaNQqQvbb+17OoW0I92qoG52axb75FhgWAAGTvyY8D/80pHIpxYlpdj
JrXj+anb0C7H0/L7a2w9NerxcNmUA2rtDS2exKOAPiRg7o5A/WInBS92TuXJrk/MMkfMiYQG1xEk
Zjh4VgVFjSSMby21ncIFwYxAW5yLXAGbHV+AmKhCp46scAaJiY+MMLEmEufcZe4xRxtdJoeI03ar
JKM5NRetloocGxqkth5Eu6uOzfeIpHa5sEUGbo5cqtPSSTEI56ZkfpeWHeMZ3n9ikpapGPIIttwb
KMya9cPpDmLdY4Z1B/I2ARjvNaxuqrrZdtiB0oDHlmviBjPRlpNKTp1fclLmmhOcA4WxA5zafDGY
Gdd88CbMOGX+pR+zCi12mPzVv7GHALc6/jMwvg4SxIs4eaaq5q+k/eFzBB6M7YqlLPumLTuDQB0y
G/LSfpwjDXoVmBxZP2Mavd6nRHcDlskJrmViNEXB9lblTXw0DLMKHjhkJaMti13i2feBDk04t5M+
O6+18dTBqIA+a+IC+MGTTNn8Ec2ihhQO4bnWtQ9rB2P/WJUUKjclbWC2gHyLm/4D5LTMWQjaDuEL
r3isyMWoWZ087BJMnTjQ6GPorRHsGw25tEkm1g4PPAxYfW2s07YIp2hs93JZ0dQP+qd5ZWXYSWxQ
Es4NAoTzNTd27Oh4wv6cEe4phkLEZZd21dIMhBwZy+n+IaRAdoRRhw294QTJhY4N4G6dI3GaDzX0
iDH2NMPKWZWvtPaM4pknF2+sW3fH/IxP7OREjwq4fG1QAdnxFksoO6Nx5dEAhFFfeo2LTAyUGjuP
bR169KWqbVbkfEJhTVTYFUGOtOCRGxhrEKouJcKLf/fJIkD315nCe6MXCGw/c7AQ3fFkXR4bp6Mt
IG3nKbMSX1aZLXSJpOJijka9xOl0RnvuG6OWGYjUuN5qSPOgW6UjbS/4PRoNGWRZghjTxx6X+Rt4
PfjEIviB6G2ltEcUENiLZuPMH/Sv7M1mKUp/IBYN6cG0poLoLAzGf8kgS/TyOK9I8vfRVbb2IUna
njjlWDYvu8z0YB2Lwqlre1C3Ir5w6IywW11mb22G/icSYNZpscDl4rP9tQxg5aT0B6xu0aeIVCQ6
ZvQ2ox+dViYjlzjH4OjyK5+n1cyLd7ym1zgE+YQ7ivBkDLPcQe5UulJi1YiUXxwRZS54isSI0+/N
PuqBpwB9BXcl4bYJVX8IkXwxnC4BqJbnPUgAyBLXGmZhxT4/cd1Wx05UCGVAcUuZwRAGZBwGoiSi
4qQu8ysFNHRkc9MdygSlkE0G83dn3NZKyM3mBmDZG/nNZqIal226dKgjxrHsb1S+NvpZ4hRHeUK3
y1bYmdcQyevIyxtRm7Ga+eWypK4lGKiE3E7qnaGLo61KHaz2JxzSv9uwm8tsROQugUEyawEs8K1z
XJ4K8J+r6qZVbLHP7i2kKex5EWaQdLD1IZxUYgZawX8q39aQLPsyFVBV8lAdwuhWK+BASzrgZzLH
7qjs+p+4yTiSvScwMvsvcUbl00KoTDK/WMH0j4ws4+403HcGjQVlI70v9b3UrNFNhxQNxkSS23Mv
8YEAdAB+xm2ni9SPQIHcsEr6lxYu1MmtoL0ksPWw5HIGti1SvRP4UO2KS095ryUZWTnTQcfemaHD
1ssdsNIJA7bjYV/ZwpkVFcFcNZNkYiApC9W6hEu8c+Q04mW70kU+ZCnMpmDQUTMCBbFP+juneFxq
KkYxSIb9VVQtS3CavyxZCYd4iDpisAwb50S5693TZ1+LSwFDoJfCu/6OfSdsWp+hmrobn1ruowUa
OV1Ex0HsNTbZPod171c6XDAYwjL0CjesaFYN7i3WFeHxpIKenzcvtvdiaXBMumgS3LRefWZDl340
WMuzpZFuvDlPhYCwmdch6eEhxHhW5IfPVaPtkSODD38kIKu9vLMJ0Hg3o44p/iKfE87aeT27hV5/
69cH5iumchfxHFSQzLpEkHW3bYSxxWeD7a8h78JIJsX3NNg32cU+E1IcktfmS/pISlYshFkDHbqA
IESZqBa8WSqDDh0G7y3AV3o5jFyDOHRJXdmRU/g+lY65ga2w9YgNxE+BJ5euCyTvZ2nSZv1mCWb6
SgYviLgKaLft5mY/aO6oMnmTzD9Lyh3F9vzlhj/pOgsYqb+Ohr12KDMy808yRGcgWo9qbCqxo/1t
4Tus2coeeiuB7+HKfnYXrXw5/lIncsrF7JFaopmmG5GJmFUzPVGBy7SkIh8IXQWaD9jPxc9a4vlK
nsY3IIa0jEJcA5mp1szyctJg4oGO9cJhe9sytw1s+QgIlLI2Ou7M1i33yUXL8rbkxwEcKmSTJw7s
cVUdi/k8PdHGUaarQAq4nGKUpy8z/2LL1gYpPlkHd7T1VDjwTpYD8zMtv6XhBEF0dNlruZ7qutTS
h11zQH8OaSBVGUpbCqCc7+0jTBma8F+9DOIgnhBNcsF3RdCHHsCj7uUeMS0rNln9tdMcG/iv98DG
nmm/lwO4j7+1HDF7KHyGlv23yT1icHHoty40VhtEjXYf4OCQJDL3REp6chJpXaR+NbhFIfR4+11u
uOJRsQEZUFlDnAqnKsUJFSWY+HSGaFoQsarp3MVMN82AKdFw3yCqClpIwSzBOKMs+bPG3CAm6mA7
9hiuPbpUiK0dW0KoPO+k6ShxpPwlz1ByFdSyRdrqN6Pk73AXnb9PAbP62e5sXaqlbyuKNkO7v3O4
Oqzt6g/6XaCztTsitfxc4q1Dk/62kwz8iOKTlADfCS1iQ1HJ+gj3RHg4M4nIp1unEiz/AaSH8BVf
7uLTG99lv3Y/uIcwLOXsoFsdnH7ErqCp8VpuSspDrHlQb4Sv84cxJ+vJ5R/A6jukn/b8i+W41BsN
iyUhx0IpVEpr07/YkJ6Y0+tQ17R67aVbtAbsXqIkyOuZzZlCJbg9A+PJTOfdMCpFMg7T0Rv6xqRw
0Frf0JiYR1UR3lmYDsFMyCxsrfXOLbbJdHXwPNkFA76ogYYQ1yLTwyOrA9aTkbB7N9AgYrqE2GfV
0LzTw2sGfL+XFNjqkEJQQfEJI0+aQrnOFj/cBxdLdTWj7wYXLbYSCvv24qS7Y4GiYmmceUmFbwhL
iFs7CB8uXA0J2ORAboyhVig3FxTjYj2IvVFMvV9aPPZtVAeQXii0KwFW81xYb57rZ1imR0GIJ7bD
/56SojgiBsh2EISgx86CYOCuV2YueMuz4IBGTiDkesuT1cXAXU8GlV+lt7RaxE4hJxEiQiWo0Mo9
cy5H91NVaEv49QThICFzIm66HS0snSXVvM1bd+zj7HqIWeRj7GpwA6cr2tzIi6buGacPYVNdbNr/
BBC0qOGRMREt14z9/st7QHJIayPtpCw2KCIZmNYixnXIo3ETjq/oBFcIvhXxtRAKMbGijobUsGeb
Nf+xxk4RBJuH53b2wG4qveqka+nLzjUXK8z9MSpx6J3RPTiKGEJLPwf9Ja3n+Guy7mRrmkJyAzVU
mLsm0uUBFVy4XOi+fIuNCq8Q0inuWepMf3Hzvyhkf6kkp7EGWsNjd5qUlk2x2oYNmdD9+MHFzBAn
JE3pZIAIwTJkZcyHd0Vr1dsdvDXsnqjq4TVDrkd//k7/9WqySb5nX2L74B8G70PUx/tJxRJ5CXey
NnDG6F5mmOhIjEEN/wJ3RL6XyUNk0ACVtlIbFzZJGoSlZ8d0ktHsqJG+EjugVNe1aNjeiDG+tkIF
NQ6P2k2agf5fyOtF24q6qHRemAejlC3tJLgnuS3UWn2JzLaNOP8EgZQKy83xfmB9cwmk5bLCfj9I
a1RZNZI6gUNkklByaYK7feregEdmOzTVNQL0g0FKNxrLzQYAzizIhmzeTMuLDSa8vyKvHBIJQbvX
VetE7pfpOCrtieL5asTbpCMPsuIWdnPAkTH+fg8KIfNb1K/zEvKmLwb52pZc2H3McW56kLl8x28F
or0zwmArRra3So7nPG1iz6Y9cKzjZ3D8ZablKHYfIalwJ+IOQ54oFQXKm7tCeGyLN7EchsGeawUd
YWi8xXWLkdbRs1bj8LWbvAsYhANIuJAAedwFW69rMbYDpmH1Z3G2eXhz4w0RuK8SBcFnxH1F+dOd
iIfKW7ugMwYH2WNXAxUaB4Fmw5Nrva7mZjSE88CjN0YAiBwgtZ6FWS/fdu2nxU8lBbKVDVWPuZnO
CZmYFhEHUplyjMTB+8TnV/l8wxZh2thNEDI+GG6SO+WmaYweqbKHCFMCrye3tpjl0KuTP+a3ILc/
t1Dwo6gFHTi0PMdGzSuQWWiQsg1/zh4J609uSukAtvWcyup8okpG/2j410jMu2zDupQ0c1ryha8d
gLEDhtirpw8arDKUkiIG4Vi0/7jevtmGLPTHKhRmI1gtnP0TNC5NOKK/Q+428hurEqvqtDfcLGUI
afuYbhrskBjWp5PCzTpOG3GRuHgFHQSaYERB+C4J+VmnpvEGR+GHoIGSRbwOj5JQFhQklSPfWhKd
bqUgDW/YoJ+gRbKU3KGuv4yXHSMARVg4tYPMdB6L1cWcAg9CLqMAYjZp+GrDV4y4AEpFwD1U0N4h
JqBbpZMp9OGsa1avm2ONqB3ZwsasYW15igToqNZzWNBmlhXp5/gnQADq+N7k9cjh5PyZsSt+zVVn
lzu/znCYqkKxdwzI6xQcP9B34GXNNUCDFuoxW0MckRUAu/LvbrY0NSZKedb8T1LXImLFE+5tjHzg
Hx/8HtM8P3lcsxDss4LtPiElvTIfcz8M1pFVaLu7SPd4X/JCzKGIc8z2Y2FgD7O/wdpChZG2+LZW
VTXezW2c2aHH1kHVIjCT1iHJEDPCnlOSqa4EinmODYtr+nlHjY648WlCO7Y6584iMoUj7XK26xFY
i6RqMIQVhpOk7qx0MLZ0NS8LFQHolaNlq9QYavqaSLccqQ+Irbl7hW8gwtflp8b3qD3AzH7bnywe
fOgYk31rt16PjteyRNoDoZIuIUkqusG/HcXcf7cnBQo2wxWdCjzN3773iGoKe8BJanITzfFm6jKX
j3T44urrZLRKEh9s68svt97+9DXVpdHHP4Nt3zLTRGY1cqo2p8dE2HyagiapfB250mbvQRM6FcOn
Pj/P5XvMa5zac9LzVTYxkjEs6wYbSmAELzzsmb23V3QvU+fxfFdpLV36Tak3Jpu2nUuukTo/YgP3
HCULR3I6U8bQLDQz+Newy6o8RqK4pLMuPGhrbKiYKQiy+n0tK/r9lrt6sg1G5T9uJsAUKyB2Xcrq
BZhmawXkdslqKWkVz5TgMU3724FDd/y/MRvP3SXh45kulW7YQI2jKqXdG0X/lYfOXthjNZYD/Ib7
KsDXlgJYu1OWqYtEHp8KZw13a2lTfze4hZZvhNd941dcH5NQE8Se4PhekN2+yp/m4QmilbYxYzBw
7njeqN+8VtHKmUqV3BYhc/SWOI4LUmu8BcPRIWIu0/xZscbc+pN0nO/Iw1WtUASfTyT5olkvRhhc
x7m2nv3nkw1qMCK/txoJNoLrTgsfcWhlKJLsFgFsImupP4S4/Owifoq3sdt4nCqV2KOL5SsJa4nS
6sPsG5EgzWrRmjgUt7LOFFzd3ozDKByyxv5uD9dNVjpw0uvOizuKmN3WkUIQrXWyF6LvOef4YBpc
B/i9NDaLWwybcdcz1E/mL4XSz2WH/NEKgrkw9eJ8VC1Yzn4C3uXqz0o1k/ib1p5DZsERdpiD5hPj
6umHKTC8QTMWEXOz2j7yfvtTyvrJdMx7oeb+LjRrqFE/vQkOoZJ8cdvsAHPY3jtTSfBvtBTb8n+2
kOA5E1ehRuxRHQoU5R+JMkPQZ9tFvM3NUPwp11Bsliuc5gCld4nSF36weR9Qvm9qhvEJPvWdyKCW
pX5ZZG0tQETmTTG0erkHag1/2Z2ZofSlyOjudz0HpWplMKoN8Uyha4Xgp4H5jJtY4ddSMPQWN9Up
yTeIKX0a7T4BddYJIFvgxoyN9UyWTDtVms32ohVB7SyGZpjVxf4zeIblA6MDpfeoOE1W1C0wAeyv
tiMX+E/H6ydeMfiyD93j4yQlX73O9VoMCIo9LDC0uzfWurQjcaknT4lbWRfvz6n+lUr+v7/HsMla
QXwm8OWHZO4psqA72LQuHypIUDHUdYh2ztT7/caC1aG2Nb1KsEvl4pCMNJFm8PWIntU/oV2ScqNs
s0PG2CjDrE0IVys2HL0FrLa2UkH179LLsjrqoFIGjmZEe31uRFdBLvpJ+666aFhYj6EkY23H6LJ9
iuFcIbfFQZRPWO88bdeOpxRqRvDKjip9E4Q5A1+vVx7dG9fuyCjyeNtOWjQ3J4kIwFwqCB/bA+j2
cmHJCdoi7+om+SVcb+xdEaEF4NVe7yFxHjvIQsW6XICuAlnXOvvqxTmist9K5W6uuDXV5+eBre0m
qwZo7gOjXACdnR0NMT8xtJHh70utIOC8FwZDT/nC6hBgckMlXTERLGfw6YeAutEGmsWzQF3Vctak
DrUYIya3C/xbosdGETkGOOxBfj/yykRmBCrBoxVLpD/lisQ1B8ZR4JD8ujeRJOCfTdxq1IpMW0p3
C+XXUG5McM/vmBq/1FXBqhpZkwSu/joKxgWFy7vdunPEKeXgyve0XAtjeGDbCFmYOij/+JnnhXQe
VM3lYez7dfUrGnFW35woQBoHPVG6fIY40zZLxJLqRRdVVmsxowUZWeqNUTYWdZL3jf0rjOO/b037
XKbZ2Th5P4+igirUD5WvWPeOdfzCXiv5EGZHJ0AJKrSy0jp1CeXmeyAMDp3QGUpxOown04PhQ/tw
aX7a6uqRHTpAP7Mg9uE3JiJXZ7l92bqtkKSUVUz0MxmeBXqWxVXdgYg4f2GL2SU8lHwqQvXILyVA
fBEzqwey4LETJIvj+OT5xLhcUr3YM3UK9X8q4WwQVE2Kb4fhAR0uOtiMOD5DueQuU0Xx4owcu55w
F3bU3h8lAx3fxlG/KTQsCqprpN7c231oQ64FKqPWnbwYXXTa6MOuRSW0XC/VogqTOSeMFTUZ0wYi
yynWY9AAe2aDvfCeIN24BsyVzTz83CdhAJEtGG8uaVCDzQvtXdpkuIJMUixW1v2Jdzuz9otg7wc3
x8Qwp62RHU6NPVYuE5aYkvwLoLrI3FIB7xE638+uuPS/+bTLvq9OvCTCW0M8pweGtdgJKGQdn21B
c+jhjBmw5L/rX+UL5JHjJM92sOz6ylIMYWRKe2xc/SsYbngu1nqnRuZTqxF5UnfIxIkXGc3FrRte
+xDAqOu6hYdgNWK2QcAvoablXjf+LaL7GcasRFzhpcmmE33JISnkBYcpSx4HbnNiQhqFbSi4xtjh
dESi1aE5N0nULtgnPec0xs8GhtSF17Ax0hUzQCnwicQAwWuviFIU9yO4mftF5OVThTHQox8BjAIc
B22XTJ468ypEBukQEwEJuQkGigXYQv7237FGuwBuvp75ZHvDx2tvtI477eFGUftOMTXoko9wW99x
VL1Nu9hXvbCh5yz/y6OmOH25wQYa2CZgrFfnOuwP2QmnAgOYhutl3Opw05Qjx1It1OkXQeMHujdr
6kO17itkMV2WgvFOAzOSL79hH6at6tgwQ3qAG1yDJt+02Bm7YTa782VPSThRSJSF+hV/swKxeTxI
1Plhw8NI79eyRiCu9EPGl/Yf41jvW2i3zshd2XxxyFjXUuZxtQeLoTUQ4sjXq1gEhHAySfcqoirH
xFP6H/84iZ3G0LFvJC1PNA5X78hzRmxIk+Xvssggjx75y6j1QJd4c6lkuxHaJwegmpA5qodp9ulv
SGMuAsRozQTi/KCwP8yZHLC/lNt7vwnoa7xQ42wHwWyNm3qL2aNPyQYFNqv7o6p1DXZ6GRxD0elK
4GaJrDZhg0PQEAoPuPQJwoQdI6pAdLl2qb76XirUuKrnSA1lIwueRPysZH8y8lkhzXePvi89Wm1e
akBLrSoXOhWHVMlcUocboExvOT+QnbFissVlfGgAUNki+ibYIIAU+kpAT+tREwEEr3dw4QhNaHdC
7F8pDrAiZi1l6V3kE12fKsMR8YFELqLOOoCT7IMXkwdB5mF6gX/4emRmyPTy1lVOTnPqe/+C8M7N
Ad6nAU3nAVKNFq5Gr0/Weds3tp/0iTTg1M0GORlFneNANIpWzkqKmtNjYx2WkNxVTlTYxTQx91K6
bi2MjXFZKMVgWYhAF48w1myO/m+WXUZh+7xiSIodeqyqZ4hJF93C8gdIYcYwHpK+DnyhpSPIMn3L
eJA0PAl8VCShD8V9gHDtsgm3kn4DapgxSBgt205P1annct5GdOMS6exu2rjoDbPJ9tBfEj0aHLGS
LdYU0593zvWgbSJP61tNzWCE7ybdez4hCMYUZzDzInXQy0PBwTRhXIxFDnfNPvJAepYOL6Sug228
R5pbDI9wzF1bgrxaoaktmiFEwam+OECFvS5p+vJeKdFI5WX9SiBqcrmKh/mh5nBlqW2M7DQrFomY
+xF4ASxNEAiYn8Ss3s0dmLcTGy+WTSuNz2l1CLulB/a5jppQpSOlqE1cYgZQc6GKNerbp1GeeuVL
47AEY/hXmfxAet2jRvt2+63QPt7k12WQnynhHmMAyZUMcZ+EIy3bzM6ZvaVl2K3zyVlMKZO3WYnR
5KkU/L1Sc4bnsHU5DaoyJTvpRndRxL1+rdTOZ11BspwhI5mVGAFIOoH3egjzvmU445tf+9Nl8XJ/
hpgfdVDZrYexPFoSJy15CuaHvIhTFORqYAKIaRpLm8AtZo6glW++ruuIiNsXFawf1OTQT05ZYXlT
Xevwj9aH6vvensOVoPJIHgK8zuXPYa58TRg0FoNDuDXHcX3jVGlw9fDAcpCvEEpiWWA/hajgkjdM
M0mJk0oKs5M+UpNhqGyrzOOIhDML1m9t0fpFc4I5TbscdJKsNZe0cY+wR7EGRksZTlVHedgZ5nOf
htaWdqmhTMcttBdV1tq5rTR12VwfsdJvkDWHEoCe9MAhdBLZaFnMn0KuQKUctv9oDGxlupq/gsWG
BfiVSrhBNWn0M5lPlP+u0l49pqGi3uZKmnyLJIOx5AdFaboprcpq4mrdir/0vjyJxbYHBZHVpDPW
7guhhHDfognA8wf5ftQ35Sl/HsiJyrnnWlHeevZk/aKwx+9nkRPQsR+Xt369Ce4QqUxCsyMsdK1t
yaH+7YNEcveE0re43yUQ8DLSTDrlZt2OMJ7CBITy/L4TpPxmKiZGIEYF7Twk2CBBeQAxy4TGkNRE
1G1vhorKqeJcUvI4JZAmPZMim3vw7WNVl9Di137Gkb7r50lbVZ3FvaqKxuhcc7DLLnlvvLsifylC
DXEdmD8oZuMKefnar64oLHgsIotABtMjxnnoOXz4eiJCtX51QAOrAVMkOmd7MYpA8eEc8l//9b62
FN7b4Kcsei1ID9HDxIEemioFpb4k3Nl4DHymZimqCvyZ/2O/cUPccxKETknddJitAnlhHDmyPgWx
8b0aPR6UsVFgr6gfKQVKIGQ3Hk6J94SflqATndtpKS/mWfd3goj5dqP1I0CjGRSps0zMsNs7WfbU
zZQ2MV2FVQjv+xmNLIwCc3l23nvBmsuuoq5QnbVM2DR6qfSJi1/7Ky/RFpR900KejGVjy6sy9/o1
wWEen3XRp8koN2qS5B9jJmHBl1dMOrSUAJVg1xg8JToc+1qsne4hCE5A5SAnnnbrfZlK/JKrGPxM
gW3qh+uVU3aVFUYqGYSwGKGV8y1hrlDyPUCHloeDZD7AD3Q1JH5TdsBCf41hsnLg0iRdT2ZjY+no
LN5PEAlH4M0DUuSUxlGXigdY55fGpvis0tBmb9H0/WX/4LHc/di5RK6DoiAd5PqUnirdaNP0cjN/
euflmj6F9T58Ly8Tc7HuZ9I/y9YaTXpCvMIwdBODMCd+wMdN1yZMiU7atb3tS/oRQu1iu7LTmq4u
UURPVe821JiYArkdt+tLTf806gLjtCU0QFZ1g3dLjHFzYcuPltr+0VC0WByLiUko/e0/ikoH3qnr
vH560x7AaNQeqpx6ACV0HxqwNCgTbUrIs2APoWYsmpIASwMDuCg9YsF8gDsERCwS6H/yDQfFMA+c
a2g/xAdi9KY6A0hB5KxyzKQMz6lI1cc8DWJ4YK7WZqlyDQW46He7rxGf3fxasx7ELFKumDvnwVV7
f9WP12HsGnQjgo/UwnmczPAlrzZ74nd4b1mv+aFmvjrPkw0cd2FC2FvtorU4hzVc6B8VXYY9M07p
zD18F+P4Em7pEMl0KAqQm8kBKjA7HwgClBBuLkse3cYlsPlzim2LK8fQOGwpmYG0tA5QYMwTCE8u
a1fW3wpPhntj5anbzy18/Bl5d4YnKov3vQmZDtkAZnr1dmXPesGjXCWFTJ1nkSdfVJHh3BwIpYCh
LNnQha5rI5pHJaAylAUtmUP4FtZztsJXQUQhWsCoS2C0am4mEdmvuFC0o3+tkfRTncCon04v8YuC
VvvVNi2EMZ1chI85O9KI10q4AvFtsgtt12E6H86cZMKRD6F8AjRZtZoSVyxVD03LXzHB2JBoTux+
JzTV8fKgdH2+VzYqzF1zj93Uy9n7Sy+sSrl+1r/cfHLUDbgelLwkYAxS5ldB55fSPI/KveIQDfkL
XrWGFQwJnYAJRmF0aCX8ZAF1hb84x7jtkS3EPQkAhKdvICQyORfzyh4X/j3Wm0S64k8Qtr93yNvy
OmlE6ySSbrFq6PS/Gk5Szizd6rW+nA7PoAW2nSRe4JDi6SVqrfdizI0ChFFyrfz3/dsF+AUi4J04
WlYr3bUDuTH6PpV4obS8XopQYL/reQbibON4EvSLqLComPTAXtNGVmbi3uNlGr7nsR+wXo/8v/PZ
0Y9gz6emQZEH6Zgt/HhV4ZX+UtHBCM4u398QzMUqgBrB8wdTO8W15u9dE4jQVFgsRep5vy8oac29
Ltbf+GrPgLtzTBhDmmsyj6RFoXrw5k5ZkHHchwmorYT0n5tXt1EIEFgPUsO6PXlVUSEpJVPAj0tj
kp0yQyNx1GbXNXZHllKG6WIPoW5OIUCu1K52XG3kRTGbs8GQh+2x+Ej8YluuW2L94ilOKhWR6fyf
MUyp8WlgeUAV+kmZx0yVI1+VDRUv10DrAvo+L40XOFEWezVHQkvX95OQIR0xh4cxVxBn4cW/xImP
FVA4OsVdq2fVk+xkJJ8SyzyhoDqzAhz/Uor8XhmklnzHp4/jpdRqGVjKQMRXW7FX91E+vgIIyrN3
K8+YHDOSZ3JZanFCTTRd8LFLt9NDTra8rmGgMFrm0dhM5wDWk2ZH6mTflfgvtwyMcFfPeucRKLRb
IIOXiz2X7Ij6ZJ3sX98TOg3gcJqIMiAoAOLEoPtHFItSQDDZh+XAQqS9UtkoKIVslZPJ9IjOTgx3
ao1sqjzpNNv4Vvs4vBDmPiSTfhZIjc+LVutv/Pjw/8arqZOYWon/cw2G+hGLPXgfrEVA03sEYwmE
hPVWzrH7k3TGowplmjO4/7hSOmt7IAhFHH+2SqqfV8r7Po7jtWW7ME3G9NlCaJD3bzTnBoayDiBp
0XEc9C7+J1M4D6DRDSrxAwqlX0anOnRFQIlYWg08lfbxBtyEGCWhubaAwK+ne4xiLdYrXBaIonOl
+qYFAHkx5uWA9qttL755FaXxLrclCvkLigiglfPRrRZ/2kThUzbKKXDnN62mJieojfISMErc7Ebj
FfS/9Q4xBBuq3KtZbB0KokgdN2d4IN+XkHtPVBLSevXtyaZBZ1ogX3QvfdxzHr8LK3fEpsDrrru0
AnnpxSqwGpw2cfTJBv7Cu9ulwkTd4rlEN1iZ7L7yggiWYyNJdwabn9cBNvcfrNFk21KrEop/+TU+
6T3yJ42Xo1T8B5cmDKNRicOsCgBoO009986o9t2ju28isB1gvKPGDH0cYfdAorQxZ6p7oqzIuyv1
yGN+d2dLXy5XsHBed+KltxviliwW4PxaOVfRMrm9FB+h6DOH1QJtzPV4g+8/OGGp4042zN0rX6dW
SnZZjPHx2ui7Qgqu5DcOrD0EI2jkklUG/XaUL9HpYryFvY1mJYLBrLct4zMOhN1qEebSwcnZJvff
vDULz42JviebunVYdey1VHRaQBIw6F71N37vo4Zk6PCslEdfH+ZeUigoOK+dV8vuFtTFhpQ7RYGm
QSTsHtg0mX9MBveJcu4GJQoGejKdtE7WTzrAenYKpzD9Kp2+Nol4+7ywg5eE3q3Nt4YkQZpqn32q
ulrW5aYOF8yGWT4LqViJdAi8zOW6eKCyVzXC2I9KJwS2LZwjc+x8JBWYhy5Ve07w+mNaZVOmOnwz
KUtMdqd/w36dcwzMKl4fQ9uOgr1qF/3eQkqG9SaxNbBp61aD0cuvPNVN2/sfECUQ3NZyQEcAEf8q
5tq1fzqcMNuY0UCwxpG9ykHylBZ40lJAvJHgkVLzBr8t9J4c7vldJX3TNsnuNKE0wPlmSZ+6t3Cm
1UGmXDx//2w5brRWrtljd0e9jPNd4yWwvWM8QiTAozU37tqMfSae+D5dV19JIJpItogrVC4M7BcN
NJtDSApJVrqXc82Mn2vU4c79QOHLTo1ItBM6CashaqbigIosAbbnq/fxu6IoBu5JQc+vMqsnUVBK
UUCgq2ZGdjfGJAhNTVOlh7fCN6IsOMLJlySyr/tOG3K/Kx9cXkazt/mgVCIIzCtfyVF+MtQE7QGC
QCq/+v+bLTqwLoHD7PmXstrncDDgvyBwsXXT4TUuyb7QJMFDJHv67ME33ga7A0M9ER7nTyhUrtYo
rI0Dv6ubSnf123dQLhwUvB7WfdpQB8dzsJpZKUiDC3zxe4N01T9jpTJCjudjkNRLdlSctD1rDQVo
X5JIyjL++dvmz+X5L81fTkH4w2xwhxdzbcVbQSax7yLWT9+RRMg/MEQj0ChJVMuNrXsqbM1HGY8G
hoJ0ZBCHXHE/bhH7bRvYr+c8MC04qSlspNG7L4lIXHRJHmAJPzvzIMinUTKkmbAuQukEuyoLcdiH
fH05zWuYOjNJTu2Fzl6YgrFZ66Zek6+/yqf9nXL6NNeHxcWQEEECkhNEKlVUnnH4QiN5qOGGm3WJ
5xNc6zAvNkALIgL5wrsFIZKmAXJ34ALC/EZBtdYbcTqUIPjLKFC3lFmMlDewLF44RkDLK9v+DQQn
xmv5PQ+DbFVxSEUkmd6w46coutYW7eAWpew7xg6Bb9+VG5TQbwV2QQRX9lvTHLgx2f1blOAH9Crk
I7gXiek9IL2gn1ih0njSITydET4Gb9d+BdKNhzD6fsnZxhXsKpt6y5WTbke9u1I5cejyz59/yYXf
xJACtjk9JGYhT1GzzlQWVSvlCLIjtQIPaICUCDYnLsVxMqby1/wNxGBLcMEXB7o53wyuaAxwSj+e
8R4qfAgwwF1wm1ED2mUH/PNId+pvrW+uOZqZkf3LVib2vRE/ouSaSYnA/Uh5crz1ZzZPygkrDHsj
zInuDAtDmyvAjMfXIY1z5lrXfBSHRt2/Js9sI6ICzgUW9c1hTLDOh1OsQ90Dnp/4wc27Op8ZGW3F
q61INUQQT4sVheEtHhx2rmD3FG02nzoXgzJKUi4fawWUnUskdd1p7kCzUtopoqFTK5VlMEi2zjQ6
UfCyeO/z2zVHbK39yhr85ltPuJ8WupxBzlxCCO8VUZwZ1fvkUu3DY3uvkFfabIs0+0FC3NaQunlH
65/+PHVml+8JsOu6Ah0FZGcN/kMSdGH+683KeVyVPKmyrjiR4DHkPXc9yV7R7EtEMC9imCeGkl9+
K9cicghFi5r7MWzz960ehOcEqwE5OUM0+VSePl1NAlZbpmltjXl2aZxouLNDEh07xuajash69ZFS
xEfdWydeLeCsct5/9rnqDN5IfDq4pjOENFwBUdebnlIqhv5pi73jwcj71PrAOYfgFtEHR9G7uHkm
U0Bvbk4x5v80nmpWTmD56x2TPrWst/jUXXYGswhlheMheUnsVpd0x59hW2UjbFRDAA/6l5sOLkkn
xEl5Sf70v9WV3LVmOoSggESdzlReCRWIFgU6mJa+yM54YoKH6Dwddt2UuQFLCBgolY2bNwBDEyhj
frpdasjNNQOsLyzLcLlK1Q6d5PPMwR1CMIR1trmlRXKXlqrE9kH1Q6LmrybwL3zjT0HU3L/I4rG5
UDk+gw9F5EJRP7DyRpYhXaHug6uPJnSCazh6uhzTjK0JOD9Pw/bDLQe5lMhUg5JDSXt6xoRKqXfu
zGK+X/FpiDyxJxZR/z2U4hpmyE/I4hNNhwmjFgvkZDRJJqe4uswY7b9FsfP1PceiZvyRvKbjO3Ik
mUZIphjenNG/kLjqT1yNdcN1JkaYwfVl84u3NXoBZZnYGqcjdCBhbawqZ572xzodx0NkrFJe71iG
p7HHYLsPVwNyoHUN9/8VrHqvZFVJ/qxjDBG7Gr0Hn07shxwT56U2XG4WC51FHBkBeQ7jtOVee/mh
SKkiTOK+5DE1VBdhrVvPT2TzTMoVR3jPYAXYcu1I9QkzpZmelmbUhWLA+jjPfZXZUPoLRelBJPD0
Afb3RTYFicxBhATGKZ5PCFRJ2kZuF79YCPfP+Uh6+ceo8GZaWb4PZGXJSpp/QrPjMrLIB2boEdbr
nNrCBoIZ9vpjDhN2D7eMT94/cbRJdjDoWS0Lj9LISih0QtgieMz+p8JP6pXSCkD8zDM6hLcC3Vqx
LET6WNPfVSmcL34Y1BzEnTb101wql3FOO7AQ3kexez3GK7byloyODwbWKDri6ngBSdaXw+HWfgkl
fJiN7w7GvgzK7BxVmnhH+Vm5IjfvpKq6XBZlZouwuI29hGIPX/QMn8KiexleZEJGBceG7HoFZ8xK
ooUDTXXSeEYE5g7M6G3YPkszpzJxntJXDnk24iHt8n5QFj4BXfmhc/Adnfmh/Kj0RoqvKkZHVR92
eQxxrAA/AMX3UN3IfZJ1TK4aEiKwXfKMb3K3PnghuOPsXlWdLWa1WtrQzxw3hMjwd/S2/G2F6hGd
xex81UtmaTkm0hQ0pn8LfyfrbbIy7hlU/F+ZRz8FgiRvKFww2RRAiQc5iaBDq/3IDoaODusXJYuq
PnRxsZcC+N76eBQrY5xsfQuSTAXod+ECQTSMNJ/g56mgPaROMD4TQjdWSxhmRzn22S+zPvZgypw2
q8fzKqQSwBmS144hVHqXV1ZXtb1SbN6QZUjk69g+lWOvs64h2UzuW2iQwuOMyLj17JakC0bVMFg7
wzP8Or/to1KVa9EZQ3GDRma2w4oAhP0WHYY45KIsrAAGKzVBnLOs1LilHA3D0khv46zFQnGkl6q+
V7+QmGU5TskZ7FJZlEwwMG//q4I83Pn2IgcukCBWsks8D3CxGvj25GjVOJOdcunqfJQOOgfe5auM
1grnu14LSKqXj7fF+bDA4mZ6qtI8V+AldlutV8sd31LpCt851T3BJ39z3o+hgqwSFr7CcuTTZIoa
KdruJPZ4iXZjUm0vC6WgG8uI6vcDXq/pt+hAguJYid7/c+/s8EuGvC30nGBDdB4uncuMIaprsLpr
tPDGa3adA17MerI0O0hdZgAWnXCwUEwVsMsTxFTwvEGwK9vciR9PwJNRp3CckKupYD7FLoCIWNQz
Qx9PhMJ8D76Q7Nee6tSO0avKoeqq83KfstjTqbv1HHox1ldkkYhj67RoRvo8P8wLkA+fpzsIje1v
5NR+AgQ7WIJGBywStUn6WfDyPmiz55n/pG9OvgauVdQCPM3gr9w/8VDLcbsL4XvjPzuWIn2ZOG0v
sBI6IU7B4YR6n5DECeaeNen47ppNAD6e5NLl66qMDSUGdNwSlUQjkilvVkFPSX1+3AOFVlfXs1zi
IWKwBVPznovsqFLeeuJiFGmnXoohPJ8bEuwpbHw82VHLXlkF8K55VOMU/Nyl1TfLtHN7ZYinLBwd
3zT30VX/LrxXTQw/4H2lFnmfx9vY3omuOHlEV3viv32x+PJkAd0l7L0FQmB24XmJefJyDqod1r/l
yG9OBMtGcnr5fPYx9H94nrTLD82G5oLc5vuAmbFGBSHPQEvo0w6vIMXnQ1UvbrQ5vn0Bdm8J+B0S
9ERbyE+s47BoiM5/nQuyrPXdO3jK0QGqTLJcSNxjSxCh0EMJKtnyOSxUywBT3jZQSpI7dSkojV36
mLl97yQzSLOgVwZ6ohXVLkCbJJ0z81mkKR2weY3WGOZ/nWG+5fzuDgHqrtmQdyMtUomksIOa/IhA
mbz0keV+5WAVB4LNSD1JTlFVosVX1KMmF9kh56HKvv/83pDc49X+sDq+HkxEhE4F3eBBShEcyGDT
uH94iKF+9KdFUyOdCsauvjyDWoet419Kfb2vKoFAg4K23eEc44+TRmxSiE5M3ya8+OoUgE1Eui3Q
Evzp7tPqg9gwfdXwAm0gEo+B9fks32zEDmuothjV8+EQc4garIlrrsLuuB2MLMq0qV5dyrFYEFaN
MVl6foqSTn7hvIlDn/yJHgqsF4a1sk8W+gmgPckOJd+uk8ZNUkOaTU5ECvdmreDWz3q5uv78B3Af
RrREVrC6QKHhOWhpDe3AO45a5+n0PhSaICZ90ti5L1MiKP7BpsB1wMBO/JuV61WyziJnczEgXvfB
LhuidpHI9r0PeQJbFwc8UIRtrC29rxXXbe3v2kOcp+OHeQl3dJJvy1Llu/xN4thCyrY6J+uCtDTw
jJNx7tb0O6ENq9G8MOYoGVCTs6zhy6DbUF8NsPlLq3bxLvYBcMBjsx0W9g0W2bclOPzCVZPuftRr
UaSZn4H0abzZsW3D+zXeFvChpKy69ipgCbRQaOOWHihneZ8RU65eRjYdONNqsRLIfrwEmEhIEV3T
AIuzjJCP71RW1WCn3HvK0ZhT0R3bYh+RW/aWcExjNlxrh50bS9PwzgrwU1d+ZGRi9fpaD37+Sodt
Kl90dWuWydhzCdlKTNWbwLCpWqsH0/PFoonlsJzUxqIjYoyVhXqHcPVUW/HPw3x9BixsUCnS1+sY
Pqxj4ou0FXPTmk+kCrE1ztxHV8N0nTPcANjIgYYevXyD27/xdoCqU4jKPxc6LUwpFg9mE19NzC7q
93ERo4dcMHIxBLT3p62hl80if9hbmFk36hDpz9KIUiCCMcgvVsgQO/3hgpVN+BNLDEHkv4YnrgyS
XjD4UcNGlWDVafzXxuwPjhB29FuHZ2t876AZi37jg+yYCwFm4rriQLlLN7y3QYlMAnV17yUGJATO
k2uWoA466dGyySPSc0bFRE+FaqEcayvxUqDT1kpfXetLaAQX+FXzurQdpw4vXRBOjNAtncTeN7n3
KEa1c6ld+LDu6jP4NFyD+Euqa/yo/LNTrFb82x3hiL+s3gekJfBDzrG3Npfgqly0RdhIDQjamRDL
JkiXrc9eShOPZ/2QbIWyW54jPoMS2HPUx/FECahCfAWsAMoGg6dZIc2I6EzpWBxB8EkjfbJDWONR
jz8I6nuJfWsI3U4uU04nsbDQ56Xrd/W4ERkHne//EC2wDoLUWcKzn2Cg+3J4Qvjv9C3MU8eQu/X+
qWRMlBiJoL612i63O4IdIondlRpIgHMINFaRCVqwrk1UQAA58Dj0Yj6Z2cGOst+fP8NGyJzPTZ3Q
cKFsXK0HwDWnmJhZILiii+rBMFmXDwXTTdYJ4v77sg6pDS6o2vrl+wHUQ6W+e7lwWdXRJbKzNjfz
PRtwZewNXfZ81pMym0vLRW2ZqARxkJi8VmyTuO0CAdGxjO1FDO0zs4Di/qgj14YSB2W3wLWXJpGd
3xlM/1xDzQrJuGArKGT4yssJaP54eCsFpZpUWiVP/WwKs7G+QyYnTXf9toSRpskfm4P286eFQ+D7
nPzac5y4ho6+bXY24aXtJ2jM+sSbneaaAjVhiIV3B0X0L7Tkg94J9ASP+Z9TI+zXQKx2bVQ0ioj0
iNYolS62YVR8iQeAdTDZP8ei0Byyo1hs4WH3ug4OLhPxZjLdOxsnVaCANX/V2s4GdzsEXyRXKI0O
IiiUSXi15Zf8/oU2O/95Mkk17I7XzkxJ39bdIwSAvbgTteAqET0x+C7QQIwTjNJt+8J/XkkqGbe5
nsh6HGKmI00GJ4LTZVhQ/qb5Jjw+TosUfeNUlBDOl956qBqywTQyxQkrKntTByioKxhpyS7bppEP
NZ1rBzV3qTWGaAvrFr4DTOLA9XD6XhB4+5gUtRSebMqhO1J/KZU2E0NpIHSPykMPLcPnfxa5D8Of
oy8PrFvb29hO6FSuXbItUBG54T4xqnr9+NaIcYClqc+iWEzlRdH7XFVnCD5R45Fkgl2lvsK16cMt
fNy6xCw5R29xWjtXL7wduzNKaSNOHYwmrlHmy47HnJA0QfElQDOEkhgOuZSbRM1cNUkIvhKR/4NF
6OwVx9EYdmGMLRxZfDCuMXkDaTcn65n2jBPRY9ec2velQuYssHz4zjOTQBwkmQvq728EMpgOoFFY
rhY/HdwVPThKQg5KepOOdk4kLVV9hg+4Kh5e6ovQ0w1MtVtXBC0KyhpbWGo56n3IZYpAuH7NHaN3
ETke9FUFPNy4kdysjp7vRYqq2OO7GBQuDeNjHb/3worbrFyIq0WUL0EMT/lugpUMgOr/atXjy2jQ
ioLq3gBtRGYbMhJ53gHjdDTdtsDg2A5D3Z1VAWGi1XyrpJ4aAu32dSqrdV4HslSS38VhMrmbfQUy
IJWmqOrf87eo/G9IOBbvhBJKGHD7rKp+LHtaCvmIQalEQpZjZaUzDDbyMobXdWcBtGAKQOGhb2rp
TVlOj+1IIYSnSsn98TYAYPXjdXtiYweI/r+rc6cUa/oOTfaiht0o2sE3+/oah2rHYdcp8ZrZpSab
Nmy1iyyxKbcRlHzP1uz1uSP9Tj/as0gz9L345Ud7X66ZvPNF1AqqnjQQSPffn88bhElahF1XR1LN
SLTtYpJY+qMEui9+U2jTgaROGXagbpnYGy26zQx/0nKWwsHPNmW463Sl/1fIYjvcU5SHkyl3QSBk
CBqKpo8Jq6KERlSHzYJ8BrmDoLA7gVA+5mbvjsQpsep1YSmzk5fPR2TC3MYW30D8daP1pvFM16zL
ILu/ceBnxGKFqP6SNZPY/NH9YLm1xHs4VB/DUJWyY5Z3yc7luqdwX+FTdCp+2I3CrBiajNO505Dg
LxGK6DSvEz8sMeXUrTxpc7E92xPpWPMRjgff0KhYEbUOkgZGa0Az/iDrgeXxZnC0UkA0t6DtH0mB
8ILO4nTChLIfEaiDZiWGS0jacpTrL4uj2YmTZhidq02xKiXMmuLLDaiEBivyyQIP3U853Pqm7+sl
+stKryNU9VT0tivmikMwa3jvoyPG86cgi5ak7gZ1w7f0oOsg9WT+ZR5sZq1woR+bwRZBpQtvGFIC
5XUWwme6+hEir1YtcgIQaRE+1EZfy4+/TtPbpq2lsFtYvZSuhfYcqnMFf8gflrvZQQirU3iX4Kq2
zpAo58r9CxfKoeoewUsHA2oIZutDKetAbiZxX+ow/VMdxfPgSOtdrbnb3zqj/mlOVUYlmZ3zwxYq
tB2huL11f1rO/jsnUaigFSEZZHgOPi8GNamnGHxWE7nEUyEPhshyF+jzrWg23FHc1Tk7TxUlbKOk
SOgfOQmfiC+T+9gLx80ptAN1BGYP7wqLdFE1OsZ9BWZCKwkXmO2CUPOr4v8GxpAvkq550H8DGRHG
axF8x3rCz1ivulFIwN2CkxtlN2QRy3uk8KlFlrdIo8p+zyOnyM1Do3gx8tY8I6JcOA6BOZIx0zVG
QiDpCjoLeCWkHHdr85n4cdofz0qe0xqrAAQc9yL37l7M2HzpgeX390J8O0jW22pTHdd4Ngz27Tg5
QwqehZvFMakS+hPIzoLykW918qVe1TNGA0flmZhXqpvJse/werR8aW+KE9scfRQbfwBxvXjnV2br
a8qnVGOXsl1jCH3WWHgaO5BeDojV6fuQLsmlVkylfb0GNaEgjL2nerPHAKYFzCSqw/7CpjF/ot5G
8/7U+POQJIoiUAHBAViedYhnqRP3JIyP2bylAuG8HRnSmtCcU7SJk/bnB24NuSjvZ/bt63tyaLVZ
pSVntRjiQq3AyGnAWLcL6t0Nfk55sd9lisTfs3oSyrLHnjEPA0XAV530ZX6LFVFb3Zzj/Gs/yumD
9XesAmvIOCegQgqdnmRRZFJaAUbDFvFjXSgDIupFwAQWBKKn8spmSeal9G//qiXcocsgJRzz9mSm
p8SQGTXxsUMN7poRQJv78M6hSPcDLWcBbs3FNY6/dXI4TOHMoNlFtEbmdlfOXJ1gek4fTyVuObZq
LE1SbxNNqtIVibXZVSVH4fl6lnAC5vtGJ/4tOPMfAccOqA3RFog+Ea5CnZ2iS6oJ0cnRR+Zkdo+L
b6f4xV4fgunxSv2LaDrePI4AKa7Iy7F2z1YdtFLzRwxBTZPBVIKc2pEooYim6GseA/RvfU5ohRGI
PYqRYkwUSNA+KQdx9mb1bcSEif+zE+zZCSLiuF555/GUx/lLIordFO4CAqDfsPebozEmUuN2TnMI
ErSYnu1MO90r+L1jbHw6sYND33MOjGdmHj8U9E8p/nLKWo96gnsaEZtiB7ds9n2rhjlLyV9X36Sx
EMPsJvcono5T9KyADi1inUAlJ3KEoueCrrNGZSpWaRNvgeUHQ8TG3ekJwOSeyYtT4mE1Llqgdcms
SKSLbN/2VuCuR/UVFTX/M7sgFSDAUyGpKlbIY857+DXzHWjSldlanA16r3ZMeqDZrNU6FpDPKgQi
nbe3JgtTD/zNCH7uUfF4fKfP5WJ8qF/z8arL5M3jSBczXPdZXLH+sWO5znG4m5au5HQKLAP3HKm1
qcDFQqUHkzThHTBm+yVuwglCNYgDZBx7M8y79nylGiY9HQWYvtjQMY6KSW906MqsPf6DDqLf2yUu
7vxNLRcqos0LNeT+LyI5+P16cdQJauQW3tRuXPRhTo+t6neG8GPdtTuugf3yomd+BPtgmOrdF+R6
K2M3Cmmjy2qyTzsHU0ITspBogbZDML+Rc+V9mBliPoK8w0zZIQCeSvl1PHGVapsVm7r+TCtgsbEU
LnPqCdG1NhWpQTJ/LjjNAbc3TpKMdQv2lYD+6qCskmD3tLce4E49gupYZH9t0EuqjkolEMQexQs=
`protect end_protected
